PK   m��V!je�  #�     cirkitFile.json�]ݏ��W��2�Mjߒ��!�!)҇݅!YR֨����]����!叵%Q���m6Hb����q�4�>N��}��/6u9_���f=��z:y���Cv�+�N���y���Zg�O����{���\&�ͻ�ͺ\7sV0����ҩ*QJ�$e&O���9V.��s6�����;�u���]��C�K�3cJ�0ee�J^&��.Q�,O�����#F֨�fh�[3��2!KcL������L]��Y8�V2����N�	t�AA��<*yV�B����H�r���0��Y��Ɩ��C��:��֨���M ϛ@�7�31(�&jl�;f�@c���c*4�C���-fh�4�2nA�<���-TUH�T��ϼr,��r��"͜YD�8����9hd�	�g<O]d֏��$/�EbTZ)ǲ��7g�5瘳�Z#�4i���*eT��L��T	�Z2�i��x� 9�GA#�V;�-���}uP���;�q��TI<v>��&f��	�z���QgT� �c��ibƎ�&@[�qs#��b��~�bd�5�XL���cQ��#F�Ů�4�XƢG�W�Q1E��1C��?0��󓠁f�ء����c���E���tJ�/6�M�L�O��ڿ	*�O�E�p�$\T��2�X��[Y\��Ő��.Y�8�.�D��uD�A/��/��/W4l4sK�� bW��ź�
Ub�^��b"ŨѢ�8Y�ÆłłŢEq^,LUaش(�J��٣�WU��M���j�PҴ(N]Ui���4�X^����ߨ�p� ���pV)�'h��]=OМ� �o���J�4���$��ř�Zh����U����`Cs��^M�V�����0����߸���Ɨ��W3��ܸʃf��%4c6� �ٯ�Յf���/4+5B3L��,��мϸNጻD�l̸�N����$ɶɚ�$Y����V�$	�� �"I�(.���!�bI�8.)��K�^N_N�_N`N�`NaN�aNbN�bA�bA��iP,hP,hP,hP,hP,hP,hP,hP,iP,���$�s����'I�\�'p����a'I�\�%p�� uD�A�u��$!`C��^<I2��$�s����$	��UY�I<�����$x.W�8I��rUY��$l�v�\Y}����5�:����mr'�t�aY����*[��|��oꢬ'w��
<���b*�0�3r��Si��K������b7�3���Cn��(�+�����`F� L�F&D1�fd)���?����ƣ�����0���.���J�aƎ���0%��;22��F%�0Cc�a�rwT�:&��:vM^A�~|<Fu�n�އٺ�_�}|��@z�x�A^ d��
�u�;Pz� �̏
�E � �� �?OAl�DX��@��U1�1���� _"�����G�8^ tN 6'p˰Q9~���QQ��z�<}��)V�5�K�L�
�Erx	���À�(�� �X �_��.v���b��}s,�ܻe�-�#˸1���D��!��cn��}v(��lO���0�Jn�8)lh�b�ʱx�X���L(� �ʶ&���q���mYv�ʒ�>���/����âX`Q,�(��~�>?��}��#2�t����!�U��e�GT3���s�"�\��aYpIw��vq�gA�Ȼ����D�u�?���G������W{�`�@3&3���ʳ��406�d������/�����v�	���Wpi8L��k�;�"�\,�a�ʄ��Qp�x�](�:�;L�m�A�]kc>�ļ���P�~�O���er:~�mH�@����p�	H	��$,d�|8�Ҡ�Z��&$ZP�Ph7�]�v��	�9��mj�M���C�"���=ڄ�=D�!C�>V�I��cB��˘!�PA Z���nx��n��u�p��OM�iF���q��}��zJ1���o�Pk�x��5������C�� W�7���3�*��A�	�b񾇍{,>�~��㞔�,)�����磢��8ȇ9���n���z�G�z�9�D��������Ө� !���8�q���/�{/�ܼ
�^��B��6��U���6f�����e�M�}���x�I�D�I�d�I�T�I�t���L���l���\�)=4��&~\�_~Z��z��z���������������������������j5��2+�MV�{��|��6m@!�6O�I=��W�Uby��(��͖s1�g�+���|UVM�z���Y���>k2�������湬�e������^�mS/׿����w�{h�N�g�]��m��	ݭ�~����}�|�q�W�wrWe�m��e��r��W�鷺��nY������.[�l������L�}}�$�i{��i_7|����gn*��Y�W3����u�k�db�f�Ul�dL�˥�%<�P�-��&[/�}@��dS/�ve{a&��ק���X֋Uy��{%�LO�2?K��Y��_Z����I�/-.��H�#y���lq򥩻�gM6�+��R,�K��^�ٙ:��N�_��<���P�^�����]�ގPi�2 ^4�����d�J�q6@�@����J!��(�P�.�����{���������'|�����ɿ���_9�ښ������7�g��n�4�zO����F�ú�sun�r�km3ouM�UU>��J)�*�sP���΋͇uO��4�$��?||���#��L8����jmf�Z�P�o��	e�s���Lp�S�E)�Y3�R?�G�QN�d�7k=Ӿg�b�F��'7&Ȩg*��m�;�f�:�{��O�Z�s��4H��r~K°���[����z�|��ŨT��ֲe`M:�,�{_j�7L��L�Q�A*�{�����0���zd�����?����"��ݲ��ͺ؅>~"ԇ�YM��TFZ.�G`�̵���Vu~��B��*�$�K\Q�ğ�,Y,/��ZH�w<�ZE���{��;k�Q0���X�{K�ǝ�t���<�ѫ�S��TJ��i�!tQ
d
���l�?�m��)ӟ�����"u~u����ة��Lq%Sq���e��e�i�X+������Yi�]t� �����6c�/��x'��v{@��E�Qr>���O����[9�޵8�`��V�i��.O���s�5ei��¥r�V�U]X��Vaޮ��Ͼ��w�c���Ψ?�/��hH�lv�=`���p�=@oܥt!���e<�I�3	ϟ(�'�[�ϳ��ߞ�6���B�Y�}��������%�P��-���S��m]6��,��
O�ɤ����x�����,&���y�\�)ڦW_?n���b��2v˪�>�L)���7:�7�u�6k�Z^&!��c�64�ܪ�m���>��ŋ'g~r�]��-UHE��m(�>Oᜨd��TRِ�d�.�Lg�.�㧇�'��K����B	XCXFXC
XF�S�w��=(B��>��\���%A@`��=@������q�h `� ݍ�h�K����6�z���0�`X�Q]�a}g�i�a���gE	2F����Q��U�27��V���IF�*b��c�%	����,I(0n��F`�%8�6�e2/6�Cu��3�s�@�����_�H��A�6�#F���p�hth���)_����ch�P��=��BO���� ��g�&�c.!��>Y��q a5�tfS��x�hTfS��i��v����*��BN�v*[���UHh�Q�.Q�@�;s1C��J	E�]8AƃpdN�x��.�]p܁T��Ѧ�v*=l�۬��T>���J��hO#o�:]���=Ĥ�N	�-����B[R@���&Z��o�+�԰�ח>�*��tq��wcSB[P��.� �_�Dt��A�Fe�����@*e���e�������J���}��&L\rMm���A>$�Hè�>���Q)=H��WPE��Sɒ��
��+�)�������ો����D:ҩK0�����A*��apx�V1R���A�E�
hk�N��J�`ƴ���qU��݄E;��	��&8عA<�Ք���ں�[�����;h��m���t��w���A<�_\k�n��:�UU�f6,��ŕz����C�saT�]��PuH��Z�}������E>�G�'���
��y�0UE��q�o(���Zt�]��&�V�辇Z��j�c�C֔�2[m'w
����e�C��e��6��4�m������PK   V��V�O.2 �' /   images/7863607e-9197-4466-b19d-a9b84c893c9f.png�UWL��,���www$��	���:�`�%@p�-���Ͽ8��V�U]��U}ѫ*VS]��Ç�J�����3���E�_;w�;ྂ�?��";��A��R���!���?�M��������F\����=��=e<l,<\�P�8��|�������������歧������WIVJ�����s��xEL����c��?|z�"��Y�O�,�Ƙ[;�����$$O�3y�2�i�V͹'���t���Z��n\1��>�|�&v�9�g���4R��O��{C���l.�)�K�aD2@���� Y�� z��s��w���E��K��� ��JB�V�o��=�ˬ��q�Gp��z������CV�a�������������?�����	�GkW_{�ili�CȂ���a�7�v�����3v�-�	�Źn��{|�C��uO��~�/j��p����
�v���di@D`,⻄)&h����M�4��������_��js�>��]����0�<_�cI�g�MhRI>�hh�d��п�n��~��)ZN�Yp�_I����3�q���CaԈ��Jq!����5�c;�؎җ���U-J��t�Ǩ��E1�j7��q����s�r���_���^$�|�^$�-�+ވLty_x|��Lb��3�*���-�{�������4+$fb�Oٿ�	t$j��G��Pђ<|eg�KS���i�繬FU<������n�sxT�DyK��PN��|#
�*�|{V��i?���"m��L�_:A�s���Ĳ�"c�x��?-�ZZ��'�I��C?$p!y�p��G�����l�W}!x�0����G���5��e�������67Tf�2��֋���:���w�t�F�*ė���rd� �!�wC��sx��J����;�!�y2C�S�F�:��l]���	/f�������,�r���#���ֿx|����J���
�v�^�^��m`�N�r������Əج[b[��z�$��tjӺ��}�7��2F?��7io��� 	�1�g����� k�:���/�XrІx�T%�G��"g�q�t ���Չ�t&SU������.Ԭ)^}�HV[�R�3��WB������P��_�"�D�����{ R�:V�Ƣ��/�+\��+a��8EFF�����	���AK�����%_!zG��>��߃rRv+�Sժ��e�u�xƻ�薄�<��Dc#�+��@�:�&3�Jʻ�����Ī�bm�
���>A�k�G��	�Y/M~߫�f�e����'ʡ���JM�O����t���$�(9fkޝ��.�;��>WIG����_=<s�'��SY�%k��M�`�4�nX��|^t'.x-�i��>�)f#�e2�q��N���2))�{�������-��>������lڤ�����zg?DYp����aC&	SCݰ���*��.}ŷ�/�6{ōc�Qk*S�dZ�)8X}HyR����!0�n��J �z�߄��{�]�D)�����t��tt�5{��?�bnD��$�/�����R�;�E���\���d*@c4Jܡ�����S����>��!�,Y��q?("�F4��J�\��2��ͱԫ̞�T	��~�f �8rT�ͤ����$7��N��D�
4�Z�x�YtT���d�7�����	ۤRaj��.O���O�N(91'����&ā5�M樘4�����C�2_50L��#�`��p�"a=}g~��q���PAf9:x���gR�_��҉�g0%�OG�23,|��[+��$L����y���{� Z�v�D����'C�9	y����7iqw�ǫO����D��/U�ƴ>QM$��SqF�4��+TR<���U�$�
kIU����;�!�B���0/�����H|����2w�����1"�q�� E(�m��)�O6$��+�|��./�7��%�����c ��RpE���m̵?⭶^�2���>1�MFu(��S��g����i�Ԓ�v`~g����,���j��@DF��rj�y��(}�a1��#������嘈�M*h%k7��̌U&-a��K��[�|�������ά(�\��'����^H��x����ј���[�a���Vi���>¤�v��_#��+g.��Rv�lB&��<�9F8����@�*���AP�N4�OCt�_D���EJ"�&{mx�R�^�_1��=�i`f~?'k���"�#I�Y�ej����u�u2u!��4�M�����F��$#;$)�K��B+ĺ��$Vti�������H�Ӗ7O�����O��j��W̔�(�b��!1~�0�.�~���=T�Sclu��(�����e��Wޮȸ(%aќU�_t�^#A�\§���\��}�$��D�n.җ�
u��I�� �-w&_GT�s+�{X�*�_��g����#�5�i�.g�4������kߌ0�
T�b��ճ[��0 � 7�M�ɡb�lJ+6��{>i?.x�1�6I�O�<�N��0Ȉ�XЇ)'�=���ɚ>���M�Ąr�10�(#1������i�`�#g:�_�EY+����KJ��{a_*�5�<$�c��j5d��
�e>;� ω��k{�z�#�v���D�0�վa��t�;*��f����eH}Q�z9��J��<��ɝ��~E��J��w��4����m[�0ĘB��&qB;�k�X��E�����`/� �����x�#�.-�\�Y�"�-��
��*�.�r���SPU��!M���ͭ�^*eH*l����~����6r�,\/�N��}��2�ph-�j����������`�a��+�'R��8�`� O,�BL�脽B*�l�$���/i�����	SK�}!��v+����Y)zn"����#oa�G�~���v�兩�#}J��}�b�����$��+Ϋ׽��7%w�����|��F�H�� R,PI����`"~M�����#xay�1;��������A�J�/�� <�J�F -��Ѵ��eg���:�R����d��\�k�v�f< ���=�
^/'�s�kS��w�ARq��� ě$x�88��7?�b0$yt��L�xJX�V}�
�i��l��P�ɛDBl�[!�{�{�m�G��0�rf�=/��Po��� _�Y"����8���Wj�P�:f�B��������"o#)���V�G^�Z��4,r����oGk����\�+W���@̏W��(��4�?"�$�,��%3����s��^��駎3F_����x�B��u:D��������L1�jH��5���I�ݗs�س��O~<ҢV�x��T�l��8p�T(&SRQ,�4��w�X����0��;���:�{qq�g�QP�N�� A�P�{ܧ�+Oc��
%�&���qo��"тas�9�\ر�c����`��{ޘ�y���eG�v�!�p.v/H�]3[��?T����쁎�Fj��V��X�1�w}E�g㷏L4�\b�c�W��5���Z��:Gw�������/����	�ܛ=��H�����]����Eb�֝K�9��Q�=����C ������JzV�2m
'�.�O1[�Z!���{�i��qaΐ��� ��3Di��g�'r�7��Yn��n��;�Q�3�.T�I��CT��os/�)����ែ�#���'��S�	sAi;^Y����2q=���Fj/4��2���S]s�?<"��y��x��d����y�f�a B�z�4"�K���	�Q�?@���_���N��4��D���u�b���}�U-�^���G�D驪����N���/,&c��nH.����:��-��P�%�~g|a@��x�h&�(�K0j�<c(2�_��kIo�����g#��{����f���L	_2��,���%���6�.>�,4H����]��{}wTy=6�����¶�$��5~"���J%��F�P*���X�5RB��U�O�w��X����w7�2�ߏ�b�0�~�i�F_2U\�w~�� �թ&��I��CKk��<�[ev���f G��ۉ�n
��A�W�,��s��Y�N�ޓ�g�]C����G��Q^.���^��� ���k7�WJ�~���v��zOW���_!*�� j���6�6�d�����I�))CÖ'��o�d:�qSr3��S�L�7"�ӟU��^,Rt�5񫊠�Ϻ*�d�R!�Ѫ��H�'�G�K�i�(�!3O�f,����kV�~M����?|�((�_��i4P=@-ն.�t�d�܎��<d�R������6zD�1!���PU٦|�u��-m��*2?�ê�bUL6,�V�`�~��!h�������a�8�_F�>��i���caN���c�Ò8���L
����-Ђ;n�wÝeM,`3zdm�=n�=�p���+��V&H��`���g���=�뚺�j�k��z�t�{���P�^a̜��8��h�j�ʔ!�x(~R*���K�2��<�N�p�S�0)���7�
_�&�އO�:Ό�^9_�Fj�f�to���V��>��s���c5��'ڊ �N��$D#R!Q�L{�&�Ɋ$3-G�;��Y}�.&P��{Bp!j��0�k	W�����k�a���iŏ�;
�</�%�X��{'���k�h;�JdE�ݳ�����$)����܅��)Aee!�GV���y&[z5id�ډ����F߀�H�b��2aym�h�I�x�I�)��;8v�ǧ����fނC�����lS���Ņ6�FF�ANe���%S��s�K�f� �*pQս�����Ґ|@:v�0��dm0�v����ΐ��rV�Qf�	)\�|kq��:���
%�g�0e$�����q�M� ���L�>�4�����6�S"7G���+A�����ǫZ2|�疭X��u4��zO^Te��{��n��d�i&�=���Y�b�*��)��I �~�(~j����aaSªBx�Md�e�礑��V=�b�;�o�������S�	�OJ1�N������� ���"�S9���/�ς&&,d��_cK֐��X3\���
j
D=3������Hb���_1H�܀�%�;�ɍ&=S�3&Rv$�$.�8j��zvě����a���|.����-8��o��8�Y���Bd��\��\�u�o������SU�H
l���dO�Ρ\.�H�|�S��b�����y��� [�s���w6�I+� i���^,iA:H~*��4�����V�Q�prS�>`�����W�NCo�����@!lg�{�8�G/sOL-����}SkEzd1�_�j,�Z�F}���bU��&���Μ��7!Gu����|��eP�J�|�J�ٸb�8��.������!�:o�࣠��}��!IQ��ޮ4N�C�|�X���h�*��H���t�K�5|����b��C2B���tnY�~3�{
y��)��}i�fC;ـ�`��9�Zx���z��Q�L��̭5a��p�� P���Z��_+�Ԃ~�9��<Q'����+I�+�TH�����F��Y� �9Vp����E&c��q`���:������n���1��lu�e�V���I�6x����@8CӘ�t��zE�/�� �����*��qo�	�V�T4�T����מ��(�O�����'�����ĭf(�ڂ�ԁ*Eo+��L1�E�;�pf����3
h�L�T�w�j~k��M=���6�z1	L��F_��Y5��$+U	��}��⑭�^�L���EJ8�G���LKS3|F�9-��d����{�D����w\��o`�qƴA?]S&6UsY���v7�R���g�KJ�:�g�4e-��PU�cbkU�zZ��,�NN��bCr�Q)��Q�űk���)½՚g��r1��`���L�x�+������H4��쀿g�3�R��>�����5�3�L]f�F2�!vPX_��$�N�����x��
�D?��1�PA�q�R�a]��c2t&7�q����:��֗`�BS��S�l����C�9�XK@
V�NH���o]�{�S�b���Ni�f�ޟդ�͈=V��xDaL��������2aEmPl�܏�Ƀ�*u�d�3,KVa�qh�O~:��;���#]B�TX�ck���������&��0� ���^��
�	)"����6OW#4�⏁��Y'IZ��.K?�m�.4��ӗ�-l�"֌���q���m��JD2H=Cv)"�\��&�i6���R8��1L�g7��+��Yr��ڴ�{�X�Κ��I����kA�L�hs9����B��	�����=d%i���:���o�Ջr��I�bך9�ީ���vv���x�˹]�)�X=px����\��<�W�3��;�ք�j�&�B�iu�8� �Q{�g��r���'Y�,_נpx��7�|�6�����V��f@B�SF7��4�c��@��D�N n`L�D���&x��yI�ګ������Hd�8Y�0��jU��@V2�����[
oY���&�1�*�G)�g��$\���ˏ����w^�d�(����+�e��a�֗�h�ݒ˰�v�2�P�®ǁ� �$���s}V���E�Ѿ���Yt��^;ou��)NZ�|OH4���7/��FK�r{6-^}"��L�7� :N�=�=n���kb}qk�(mRNFT�}+2�=~��*�_�f�r;
���T��::�~������H�g�����1�(~����L�`�L��`�) Gͦ�4x����a��b�2 A4-�Ew�F>^A�y��z���\�����5A�Z�@U"��� sF�Jp�DƯ�#~�\�?��ҋĹa���P�b���Q��S�>­P6���nR{�����Rc��71��8�4>���ju�4ɊuB��3�w*���+o�'����Y[)f��i��[h�AW� r0���	�5(�G1�W���mF�$���$0j�G�p!�U���13r��+]�c��'f��5BX�k!GС��K�>��vp�����u#��[�US�ь0h,���C@>���{fp�G<��#�Oi��
��e)N�k]�$�ߋ
�;�4GB/%�P�h��o��'��}'[P^�%�+J=I�Z�j�(|�iY�}vX�ZO�jV,	���M1��R�� �J�Ӱ��K�%�� �l"�Ҥ����	���I���@�X�8h�1Q�8��<smP�'�1�FA~0����d!̺S������/v.���@K�E��l
.���=P|�� nt�)Y�3�#X�Z�V0�l�Va`fj�J�j�
2$�(~�&.DY�W_O`�:c����9L2�'윎�R����� ��g����h�|�6���9�ɕNnΕ%߹9��GMN�;��u��]c�w%�]4[M=$��"J�	/xOP7����E'���TomN��w�\"ˤBڼ�k]�9�O�����!qY���}�H����TD����{����[���qh��4CY',3��[Į*��u
#�V���F�8��c��\y�B�н*��q�(��������ƯM7�T�I6໡�T1��yT�Q-d��x�.�zR ��
����:&�GU_#"'~�l�R��*Z��N&n��F�P�֜vXB�S�R�ؓįۘ1���3�98j7�q���s8��mł��QE�+��U��t q?2���ڼ�qsN���8h;�{öµXngC!}G)��C�~O�M�P��:�x��1T�Z�I�6Ə$�l�6��O6��;��D�>����e$Ad�Q���^븈�^%���J��~A�+q�ڃQ_���`��_�\V[��D�̩N16�ڃr�vK��w�-��Q�j��K޶�B���եc��	�e��xP�t��#6e�(�Y4��d%��(��޳��nyr�~��/��v�Pt<e�ԈS�p��&2�y�lT�+'X���;݄�NyǙJ��;�3�Uۜ|ud^4.�v�4ڔd`0C�9����/\tv�s�� �Z'[)#�uO9q�Ԟ�yᏬ�$�~a묲�}��H�]ބXU[�1��b-U�0�[����ۘ�y����:���[�=&S\��0�Eo�{��'�ty���.��&��J����}j4rW��ʳK�P�e��Mh��>*��m
�O�UW�֐����^��zM2`��z��@�m���h�y�UQh�P]�[Z���A��N��~�J�A��UȨ �<�6:�����J����������u��ܫ����H�Y��{_�%�By{�(s�
0ɛ
A�Zs�'�m�Y~�w|z"|%e����%���N~�tHeX�O�������(�9��K���!�A�5��G~��fJr;�/JK�1����e���RG����	��nk��{�S�T�U$n�YdG�c�����
a���>�>b��S��E�\��~�s��F�(��0�a$͚N�� �����\U"�!��K�>��0�F"ȝ)��z����NiYi�ESʄ
��OO��iN,n�2����ۗ���S��#=]^� F\9�p��I���i+I6ߕ������� H��-��t-M��L�v��h�o
��F�Y���^K��Z�R����4��h��Y�B�!
�F5��*�rlH��nU.����-VE5��6���n�	P�������`@X^ф�-��������"P	������	�y�7e�<Jcŋ�vS����6��V$Ȏ@�ԛ����O8���x��b_|��mb)Iu8�8O+���S
N�UM�2�Z��lr�uHY�*U�<|����̳sc���=����ٓT*4�* ��i���im�I���9m�p��8���W�xe6��G4$��"j�د@:��&k�H�&צ�;����j ��������W��@P�aA9��i%�#��&O�=n̪�Rͤ��������h� ��)uQ�w�����C�}�-�5���6��g�X����J:��׃�8{"�1�d�]�K�?�;�-���o@]xW�Ln�R��ݜ��L�ҋ7�in*�%#p>@�#�3V����U�T^�+���E�
�ҧLt������϶t>��<�ʜh�|�x��i�_�%R�*H��E��S�J��m��+B�+�I`��T�VuG���J!�������p��v\~E�q���qw�Cr�����zf�l�Ԧ��p�}��}�x(�q��eeq���}� �%��
 �����Q�ZRe�J���-�Κ@��L̺:�"��O$)w+Qǥj �ޗ��L��rG�I���^��ή�&t}��]F�裲��L���І�p��Qfd�����o����E눟έ�d�|o[-����(ǀ��"D��j�>R:�Y�� {>�3���úr�)���w�7�n!�dolcF��4(ե����G�ꛮ�I�����O�i/�KBT$z�8��!ć7O��ia�d"@v�_�����瀩[��92��;}L0�a�=��t���~��Y��#Y�.ͅ�_�[>ݫ�]�bk���[-����y���x�P�XS���QXD�)Sə�!��u�p�w	"qV@V�K:8Ӳ�k�p�$mS��}���h��mi�O�Ot:�z|~EH�T�w�-�N���x鬛	��i�z�Ƈ+Ir�����J���Sn���U�a� �8'ɩ�CbV�V	��=>o��������<*h8#*U�C!�y>+8 痠
	��a/y�'!߱!����b!(=�/������JP�)���w��B��)9r�ϒ���6eۊܹ'\�B;���i8v��S�}�_~��'<B�X�gH�؛��)6k�9��|:)�Y; ����n���Bq�5�ݐ��T_����!qS2M�8�D�g��7��=?���RM���`�ή:�"'��LZ��O���iNT
�գr^���M�2�I9%�ړj�t�"�Ϙֹ��`�j7��u�7�\!Z�GamO=�!a��GHռQ��r�=͎K�݁���g�Se���̀q)��aʎe�w>��|Xq� �[2��a��|��C�:����{��ƂR3���ls�V��u�Vո�]W��{���.[�����v���`Z����/G��Ù/����ӻ ��F��U$P�q�
店*���Ò?q�^$Y�CޢH�7[x�o$D�R�h���mI=�l�@�<���Og):Q��q��f66���r���b�e�y}J�{J�ɦW׉��ڽ=��5/tj��ь �x��k��ס�V/�>�X�^�����Mb"}O4^�+�DK;x�>)��\���i��!���`HP����!��DQ\ǌq���	މY�V(��O���k`5xQ?�ﱭ�ǫl��.��/�07��b�nN]ؿp
�('~���������j��R-�`C�rguwN����4�a�ke����l=��c�"k5,7���f<j���G��T��ɀ+����V���Q���7�t�L���x��#N$��c��%����C|y�]A�]t��$�	z��HX�x��:&7_M'!����iG�7����#!L �5;���v�#$��}'��1Dp ț"~���̽��h���&��q���f� �W�aj�t���F�H�);٘�~�p��"��-k��5�r�Y�t��h��K�-���i̜K�R��`�+)�e-�}ҙK��1�B �u9�vxa{�0�GǙ�ܰ~�[��-4$��U�>�!ʚh��SĖ:��e��W�M�?w�����}S�I�HdzS����Iӡv�I��ڏZ�U퐧3�^x��9�׮��i�M,�.�x%y�NZ�'�9��9KKo@ި>Jf��.���X6p��O}eM��qG#6���*�-!k�Њ��E[�j�_�%7��k���	>1�e����SfiH+�=��j��/�V?f�a 5*uq�%��>Tp3)T���z)2f��­/�p�KsMsǮQDB�LP�&�O}WjK��F2�	̂/&�8̳��7��C_���?�;{o�'���;R�4�{��Cj���,_��/�ŇM���3*�x�Tc�b3"�l�$[^�բ��cuM�^FNgg��������g&kݹ�4�;����ƺ���W���r4F��fڣ�˄��T�y`�!��S���"��
p�Pk��h��q�NYy-�:�;d��-���i��/�8��T
�)� ��!�#�X�,�d�0?�����`CI�a�<��W�-u#���<�%�r��b-pCq����c�i(@���;�����D�}gÄJ�u���71Gߜ���b2�.����m�m卬�wO���yLW����t�4�
p�x3�1ϟ�B�m��!��u���:,�n29�ŝ�è,ՌR ���w��x�pP|��J)P�p����hͧ��â'gt0������+���S&�p�$���x��� ��*��E�~��G��g�}$ያ2F�ִ�����~$��{�p���*��r�s�����F�������0+6a��R�p��Y����F�<��iV���O��C���˰��P���(�<�]��Իw�hLۭ)�娪�d����LWL#3�EyS�8A^Vqy��-i �����ƻ]J�8�/c�-e@�%`l�tVs�b��Xي�^r@���Fg�@J�j��/ϟ.���[;iqY*�-���\��˟H�ᕆ�(V�?§Y���qK1��
)E�!7�ح�d^�w�o���L��o�O�Y�xcK��g�n��݊�q��E�;,���H~a����� ��XkK�C4�v�ussܒO,q�OǢ͛`�͜��N^�I��BR�j�}ߨ&���Q ��}��?d6�
Fm���r�y�g7�*���H�cԘ��Uʆi����z�s���3������-���il��Z�Y���jc"���n^ZkNNY����V?g<�d��a`��,�_�}��5+��{h�{[Z)0�B|�s���I���J@.���!��1��TB�i��m��l��+�W��A`�o�=oȓ1'��W^�^�d��{Q24S�{�ʆi� )�"K�s>����5�g��L[��WB�%���f��1�b�.��K�3jҺ~���S�jž;�Ww1��W�y�K{4儨��|6��SE�����"ϊ�գ��ey����f��e�G*D5�ɧ�������>WC=vV�;�m[R�Ҵ
R�Mv�ǟ �z�����p�ȝ�?�߮�b��i��B�x}z����u����mҦ�XBe�<��h͍
4�euҊ5�O������J���A�#h�\(^�/����Ќ��ucY+�Q�;?�O"봿������+���B���-�v�ɬ�U�-q���L�5��o��
���s�dO���hK l��,�Ђ\�*7��VL���¹�٭J�0�a1�0Wd�{�7�{4ljQ�±4���"��7KV_�Є��]��+�uoDu���f/;wICN�}�~�%yS�n���=����+�7�-o��Av���I��͝H8�W(���#��=D���
i���7؟6���h�O]��� ���kbgE-W)�'[D������F��'�a�̳��׼CUs/{u(��.�H; �©�W^a�ޓ%ųY#�G�s�#����V�������8���S�v��p�f�t#S"�kԄ�1�|b����F�Q���@*w�̯zRG�%����-i�/��v�x�B��I"��H�N_w�PzM0�]��E�x�t�5C�Bl����������d}�<^��5����/>���U�t�O�%F����.z���p۷�@�jd���?3��)Qƙ��N5F��m;(o����Cw�\OU�V]G����QO��Q���O<l�KG#2~@1�����ѭ5�+��A�4?ޓY�n����W$�}!�,�E��Ep�\^�������7�=����3���~���G���_�����C)wi$뙓9t�}>&cU��Ik�~���Є6��zek2��]�I�*S_�������qG�����
�\�Gi�x�����j�� ����/����4�gjHbIm2�B�u��,�h�5�R�2p4W�˷���p<�*��]�qd�����W�m�%�E����p�*qÞ�X��k��dQ1���6�0�(PI���;t�t��9��r�z��Q�8�e�M%kWHZ�؆�v�p�7������|��3��p�Ʋ\16М�=XY]+���U/KDS��/�t�/��Un�1g�j��κ�/�����T��L��x��)���]��**?1����Ԥ�{��P�-�oyk'��>:��X�����C�2��WB�dU�j,�S���3�VR+?`8XT��W�0<��V�#���#�1��,`da>�8K�G��r�t�ޏ��G�cH/���w�S�S 5� �W�/$zr�X�Ab�� Yt��V�}�ME�����f��P�tСP��*GoSo봥�+��_7�s�0����������9�?��$��n��H��d�imf44u&�X`&�}�l�sJ��Q��xT��2%��Q�4?{}YԆ�@AL���ӻ���퇭�[�7��a]��	=�Y�]���s�&����6�Y-X#l��
�?�  R����rf�>�I�#��N)�%��*�2:n��ҝ�~H��^�-����К��H�4�J[3�O�z8Ep���Jż���K)Zb��d�G�6�O�D�_�w�������5t�|���#��E~��ᘉ�𿫌!��H'߃9�	V�mؼ���Au�I�:�}��p8�u��J�܉ZeD��b�{�I���[��4wԈc�v��m�J�������u�`�i��:��6����p����Q��~�g���H���'[�6etK@~v�z+O�:��O���@	��}�x؅�/�N��I���[�֍�Aܼ^�O�b}��ӠPCß	zmɀ��h������3�I��v��Ko�_��o>_^k/�Gj����/8�2Q2��nXr�H��$O��H;��Xb�QmB�j��<Ñ��{������NsC�E�_����ch+����
�0�O�'�56wOS�,�*j�@�]`��l����_� C�iDA��v=����j~1[����e���Q�l�������(<�'̅�,B΂r�b��sSh�Ï-�/�_���k����k-犙�W?�M'��������߻J�>�'����S�����I<Mx��׼�7��~#+�'ӳ�� ����_x�/U�ե�t(���iqX�Y�ę��� h����^����Q�O{ϴ�N�PW����^�(▼rIL?����2����ϗ�!���/�){��.V��
}ʘ��cä-�-3	Zr|�;�}yH��]�\0�ykZ��zn�l���#�F�JSi����٠ ST��@z���Ћ���K���[Č"��|�:��A<��a�jY�<�6�S���Cz�%uh���5o�E��`K��y�s��ϰ�?i@��Ҳۻj�vA�a���xB_���А����ᦧ�4K.;�e.Ƴ@�S�� �5Q�Wb����o�g��e՝e�)s��s�����l�Ǽ� 4e_u������H��cG��������R�W)��޹�V㔜!���������WD��P�������[���,Gګ9fCE;cz��F���[���B��.~�t�KS����Ǉ����Q�#?��ؼ�st�-�?����u*���!���n`� �")t�����B�+}�R,�^��Bցz�����MS*k�����H���'G�O�j*�[�5dED�(Q��)�ޔ��yĊHo�b?��^2���yҘ5�`�
@/�4�\@6B��YM�v���yr�b�q�D������y� ��O���ϡ|�s|�q�J#���\����V@�N����� D�s7'�iu�׷u�YU��.Q��O��wc@��Nc+���6n]��M�+61�m�&�3^t�0f�;1csG�G�R��J��.�؎�D*ѯ��DN>��lo��l���8>3���鯦��
I��3?������MkΟ�?�ѧ.?#�-�؉���u\��4��,q��{����չ�'I"�pO������ͦ��3>��V��]�'ۚO��z�<��i�|�~�g�Z3�P�
Z^��-w;jh��X
���w�-�q��b0l�!�e��9>lI��Z���^�\wN�ތ��zb$�gE���|K�{�g.K%�����p9���<�qx�@Wy`�y��_#�yrNljo�Nw!A���i���_�ƪo�%c�6$ɯ	>q��Z̏^��͑C'�HƊ���_|��
�8�l��-~���ڟ�du\2��V�����t��0iӜ��B%�duS1\Q��ċ��מ]�
e0�*t���3S>j��+F���8�8Ů�֪-Z������[���&��9<?s��ą���T�����u���b�䋝���o�7ӻ7u��f�؄?��) ^=`�p�=eQ��PH>�a����G���,�a���3��U���?P�|��Ȫ������PR,�sө�ǿ����R���4C�տki�����A0���aq��'�ܚ�Az�@!Щ%I���(%�9:� vr��M�{�S�`�4-z�1�v�z9@���h1h�cb;�N49�3GQ:lg � �:~vd�#_�����&�ߋ��7��2��Ϧ�$u݁HYP�����W@G-�u��<���=1�������p�I�[0<��O;�ƲX=�	���}�MHg5�e��!���Vo�'�B���� �S~^�~�"�$��=K^�u�W��3���Ƈ��r����~���F�|�<IwN��q�T�ǎ��z�j�����qJM��u�dQKա�1���ׇi�TgE��O0��يiK�p_�1}fۆn�o�^�<<�k���$kM~]�����^���1#��O��ʔ�|� �s����[`&��}�j�e���O&S�:����T��W;���
���G�t�fӧۊ�"�����'׫ɐG���$t�aB�gVM��ż��y�t/��W�Ľ�����p�yP~���j��~�q���]?����f���s��5z$ɺ���_�8\�R�#��]u�߁�����q.'z�?������0ؽu1X1Q_�9"�z�W��R�9_�O��ZY�O�^ᔅ�O��v����� 0ʚ�r�[h���듘
%ⴏ�+_��b7T�>�9 �K�'}�4���	8K�7%�W��\V`)%^��+{p��5ξ,�a���Ô�D�ŵ�6U����g��n��o2�4+%F�2��ž[��4o��Qu��NFu�G��G+�#��YWe�!Q�_�m���͆�&C!/9��w̠�8_6��]� @��[�}�ΝY��+Wq��Y�:}�ۨR.�H/m�8Ү��R��C��t��p�8��L��$M�.�Y	���R�T_���)Օ���Zc�v�7*���M½�7��/:k�YY�u,���vo�W�)��O�&x�?8��l#��C?rS�x��T�-W)��K�u������uY�;L=籠��;x~�����������4����������w�~��/}�U\�v�m���Tnw70�
��k/��~�4�X���G�Ο�	��=�,Μ#���yg�v;��)������,��Y��8�~��V?]�[g�ѽ��"w�E�ֿD�$�ͮ��{��2�=L�-2�a��r�����
4���:F��3Z�E*��e�b����fjզj���D����C[�\�|���$��5I��h혔o�-K���rG
���4X!��rT���%Ӭ��t_��u���>�O}�,�9�w����:V�R�f�sL��>5��f��<7����K7�B�0��^;�7�ˤP����P�s���G7�H^8��4�$�biM/-dF�̙<^�!���h��j�+��7�ɚ�uZC$.&ˑ��QS��K�����vZ��w���[o��fc�3<u�>�ڧ�	j�3s4��x͎����0�A0���/-���kx��q��+E�4��m$ww���(�'�H�@�Qȸz=���Y�����8[㵕���9��{p��QG��?f]��i��"���B˥�Leqi����Eާp����t�VΙR���n��C�I����Y��AK�i<w~_�V�W.j��Je/T�8S���-c�o��8�2x����b�
 �cǼ\�c��j�i�L�
V�[����h	�f�8_� �r�8>���d	^�r;Ȳ�j�o��m��n�z��;��%*{Л')L-Nc��T������Շ�ȳLgϟ��TV������W/�\*ڬ��^�����Ӻ98����x���������"��vsZ�:��H�2���0�B�tlѵ��n|���q��_���^�7!G�dq�
F�g�IFII����m)1��x�#�4��Tȋ�4�*�CP�I�їrD��:8D:7����x� Қ��9ҕD�!y��Σ���>5�bC��IsmT��m?6x� <�����zQ�T_�&�yp��ڀp!k^��k}��D=��
�Pg���`u������괠�8����sKx���X9�L^��g32�Qac�M��{����͛�s��`qq�.]����Q)Q�-�X���v�L�ȳj9�-��w���c���6se�f����A�o����ya<!��]4Q|�K11	t����P��5=��u}��
@(����8����,R�r*��LvMD�j{k��/����V<�8lo�Ism\��,c~q��
�RIx���Q=����4��+3�?{	W�?���Z��L���3~��F����7����lSs�(�9��s�0�x��4��>��)���̡�a���NVC]G����t�t�G@��Ɩ��!w�yX�PBaB8������|/�D�zf9���g�b3Pɍ=P0��p,������M�(C]��1�&ݳ=���^/z�&6�F���Zk3m
N���k��,�l$��1)���<�gWP(O����}���(/���������A�c�E|��O�����79�ui<��,C���6��&��c�I*��1�x����\Jc;�+��`ä)�Z#�Nd�S�O�ү$L��u��A�N��Me9k!s�֑V���e4�3����݇{��kx���y�u�}�}�o�y��Vc:7��3�`WF��B.��ssd8TL��<`�ޥ�np�j2��U��qӽ1�d�� ����]�8@g2䆂B�T,�C��A�Z��L�q =�/����60��w�O`��|n�D;�6n��b�ZÀ��2�F�J�>��e�У =�8�u����H{~�~�߹U��l	�_�F�VQ�8��1=�Fk�A{�E�p��2��tF9���O�P��s��H���w�����f�E��]�GM�P%��Z(��9�,�P*g��+���z<�ޜ�X��7�a����.v2-���r@�P�|åe�X�]��l[X]_�-v����-|��{�����������s��D%D��K��V.0�����.���-��Λ��@3`�(n�=�M��LQ����:�v� ��K�z)���D���f[�'%Q��2v�����}���[����`�a�;�H���{�!�y������.�˻��o!q�mZ�w) ۖ�����"��I�7�,6����j�<�jG8d���[���a9�����@�L�J+��v�R�Ol�!�~����l�G��v�4�f��VJ�^�GC�7�ɧ��	nrӚ/
C�i`��FLK���g&�z-�;������?����w��T���V.��.�>|���Qs�i*>5l�~y��j�1�}�C���=v��q��9\�p�}�b��XzY�l�*[�};M��;�+��Qϱ~��P����<�����S}���9���x��Ɗ�S�ba�.(�A�&^�e��#J[�� K������k��=̻��'ҳ��A�D��Y��!�V$��`�xa�����p��M���'�9���Ѵa*�(/�'�����&����6���������KSxza�m�ƀF\�2D�������fmߔ�e��ﾏ�o=@�8�O�����,�]kU)gl��yNk(I)�b��֎���5갸�n�BT����y���8����M��a
����.�ĦLt���J�)=lC�xb�Ռ%�>�����H�����֑�P	ўiw�b�`�h/e_�"え���x�Ͳ�2���k�I�r���ű-/覽��&�ʮ�R���l8�@;��������-���~����_��?�������)���\8{+��ųx�ʔv�X��i�Юn�����w�}[�&�y��2*�%�c��a�6��f�5&J�b�,�m;���T���fD�v����/,/��v���Z����d�F�^g��-��iO���x�gm�o��o���=
L
�9f��ln��������x��iZL�%�S8?]������XrX��lKK�)�򸷶�?��O���:�d�ls��!���|��;Bܩ���aɱz�R!�>57�!;Пn��kc촩�z��p�-'��<���6�������v�#l��ɥ���qk����m����;-l�ڸ�u�������ק����5p�
L��3�|���?����F?�jb��@�X�*i۵&�P�-,e�~��?�u�VvW�ث�ݝm�N�x���^������w��P���Eܪ�Z�ЍB��G��� �� ��G��Jl��T
-�L�{�*�aoz�C��{�����n�����UrXȥ�s��޹c�cqi^ˮL�������.���q��jY*��T�������C|鋿�g�}�����c��*�9����IZ��t�M��1���x��aPT�%t)�ۙB��%���=�Y��ZZ�N��!�C�
�kX޿��8O'}�f{���#G��r�<���R{�#Z��i��C��|����g�x�R�JA���H����5�3u\J�_��rt��������K�I�PݮK\� _?�1�n����C�;ڼ�f
S���"ւtdX7[���)�)��F�H�sP�eI��NA�E���Ϡ�2�n�LEn��!��>^}�\�5��߭Uqk?x����f�M�B��>��pm;G���U�֯�:�{�y�O��;�g�|o�����Y�f+Wh�P���Jo
ږU*��!48P�јb}��6i����4��I[��6�E����5 e�`�f�%������E�u����,�ZJ�!�<U��0�v�3������Y�W��,��sZ+�2c���eP�ŀn��e��L[F�������[{�>x�������?�,^~�e,,����m����Ɵ=l�~�S$��o��3KT|;G�������-\9�{�S�[^F����o�?����P���=�P6OCI��Ќ՗=0ӎXYҝ�dհ�0�#=���My"�=���1͑��|����~C�˃��4�xV#k,Hu���Hot�X��:2G38�x?��������8�e�W�f�31��3���Mx��B�ަ��Hr<̰}��f���޸�}�XS��)��6ն'���,�T���1����-=x���۸zy�|�E\\9��Ƿ��c|�;�p�G�cg���b������a���>�^x�e�YZ4���]ÿ��*~\-�M�HT��Ar��i;��OC�I��P�3�9T(K���ٯ �ڔ����^�u�E�K+Xϙ� �Ne��Gg�e����xCZ;������)��SHe�ݟl��hAmf9�\�j�X��#Z�zӯ���[x��z��.����u�ׇ�����/?��nR;�V(Lحٰ֧�ƨ@�A;d'h=߫���3P�&#7�i�`ZV�8lep���a���nG�a�����$�zۈ�������A��Ao�Sy����.�gg�G��-��dp��p0찼�Tv�x� ؠ"�O%�ݭ.>�Mb�D+C��Ҡ��UH���2X���>Кgg)����O�el�ئ�Y�B���c��2�;�s��v���>���tUO�8xK %���X�BA�4=�E������%�d��:�Gb�Q˞`;$f�������{Th�@���;Ђ��0]��ų�k������w�P�����"�,���Z5�I��l��.i4?;��^�*�Kx���{�.�Y��3�q �,�}�X��JJ����:x-����0�дR�ϲ��O�����#|��^=_�]G��D�3�2��'�����WpU�d�Ne���(���!��y��/�|��^���Z�F����������>�����՝>|c%Z���9��ksxf.��Q�t��]<��?��y|��s�%C>���@��t���!��>�$�(S��Y�N����{x:������:F�챁����&h��3?�~F��k^R@&8�Q@�V���!��l�q3S9����(V*�mtA��w8��x����3Kl�v��DsgsTtϞ)��3�v��r������߽���,F��H��q>ǁ)�D�|E:�Y�Q9K#�6
�3E�C'�c��GT��8����̥LF�v�)M��c��n�mt������-6�b�cȟ�M�Q�'�9�N�|���!�ֵ��G��5����m͌�(Kmp6���mDL%�����$Hh�upx���!?�b��ؕ���^���8����．��m�ʬ`|�y�:��{�1O���:���C���"����+�MU��v��?x�ܨ�|����A��F�P��4�m�G��@l�@����SS���v�)��t����+Yp�C^[��-��<�F?F�*Q��:��Y��2���1˕:l���={|��TY
}>��#MB+1�P �i��K%�ut�QkҶ��i!=��k�4�u�)-Y`<��e�lW- ��ͦi'����&�[�x��Η��߿�1����Y,.^Ʒ�����]�`��F�S��,3��9B�}�qc�2�y��gp�<����_|�����/"�p���8���2�{ѵ�rka�s���`�r/*�*��v^tbF�mQ��Esw����ֻ��W�i݌4���Ju2���6�UT�S������-`㰍?}s���p����Wp��2�T*V�����-4���>n��b}o�^r�����=�3ƻU�\x��F�l����/a{�Y����R�1l�a���)v mO�G�ޠRӡŠ'�z��h�A��B�1Ľ�6��38�^~@�lPI;d�Xc��{u����pH��h0�6��~M�.�G�>�W�xH%��A'���Il�ʶ٤�(L����z��<zؠ��LdP�&����˖l�����0�#v��z�
U�y�QO�b�U���Z��Z����-*�=�Y�L��d��Qa����uַo_�o����hq	ɥ3���n�c�O�rE`j���"Z�$�������R�}�i�/RHS�������P�֨ 4%dS,;����-��"�4
�9L/\@���on�_�yow
�^zC�FWSߔ)ڞ��&=��俺��	MI8��=B��Y���p���f��u�ï\�o�Zr�h�}l�Fx��4~�����m��6�ͣ:�)����?�[���g�0]��.���ݦm�;/-���|s�8ܯ���=�6�sY���>����˘�*��k����6>w}�U*(T������<��a����<^<?E������p��J�VOՍ��`|�$��-$�i5�BZ�z��l@#�k�ʶ�����D������]m@�F�XD9�u_����ѽ��bu8�Aa���c��1��x�xM�����p�����U��[M�]��.��q�V8V��҄���H�')'�-di���8�àZC�ƙ����AQ	���]��*k�O<4(Z��+
l�^�������8�����mAa�)��fUx6e���<C~����K����5
cA�!
��(O6��lxc�y6Y�T���lF��D��M�����HnѠit�1m�C_�]��ipM-����e�q���o������6�eZ�}c�B�����[{��i~��f;�JxXm���m������u��.bLe:~�NoV���!TM��uTS�$��*'����x�Џ	�U�A�P��6�5����a���3�C)��҅�����춉1��0�B�z�t����[�G�ZKy�J��-�&��+_�1bO/v(������>R��q�4L(�m�A:����¶��LN�_3QM(�c3�a�g�(̡1,�(��X����s8w�y��e������=��,���4Ҕ�Z��a�]�8���:�j,�R�N���8���߭⟿���esh����fi�j�sT�؎ч�5Ǘ�Sx���B.#��P�����o2��X���#�b[�z�{Ƈ:�������-��ۛhv�l��lz�L0�n.�%�h.���m�\]��L瞽��Q�w�`�����S��/`i��t���n�~`;^�)����1-�J��|f2��,;sq�T������F�k6��Ѧm,�@oI-P��~CZ��������V;=SWa����>�Uv���؇�I(�z���b�##�_I�J�fS@'�a��Y���Ndl	h��&:�%STX	h�SJ����@a�L�+�� �5��ɞ��?�*{��P%�����x��,�2l��ήm יa:�إ�.�l	���1���Ņ)�K�33;ꣲ����f��mW?@f�>f2)�\��ċh����"w�:T&��=��G��3>�F�`�Jl;-lR�4�it*s�/^��ʕ<ͼ����h"�rP��'�o;q�z$4`X�ن�L3����>8�ǹ�����KK���e쬮�TؾO���`�](�����������Gx}8�����7_�����I��G���{|���|�Ro���|o~��ZrOQ����
>y!�{��߹����*��W��|�
���p��?�������s�� ���.��%M���?���汳�4�O]a[g��̌��,~���#^ hV�>C"��/K�WL�Nkb
E=�p��4c�g�"�t����ϥ�6�e��і-eУ5ީ3lj�@�q�d���{�3<�CV�=�G��خ��:�
��k�_'�0}�C�o�i�P���&��GHo�P��_%鶞03�@��<����U���}*�l�.Ӵub"��a����0�ʺyG�C<b����$���|��$��E��AO~�u�0h����f���H���x2���_
=BR$���˼NjA�6�u���:2��b�z��,� ��� X�xY�|¶jI���r�ߪ��F��6\�t*Yd�%���=mHc��|����E1?��|��P[T,�����}{$��>�:i�w*Zl%�'�.A	]([M����S0��O�Z���mka�'��lqEo�+]�E]�m��Ӕݬ?�~�����Z��:��j�)O�,��>r�����9�~�v��7?���E�/}�S���)�2H�|d�������.ǯC�TR�.�C��5#�,2'�3Ŷ�r�u�&ưu��oڷj�e[oݠ���s+�X:�4�4�W��:?o��}*N}S���%z(2�<w��0���?O��
���A;��z���4���ؖ4�����7K��J��)�����-ٺ��d�a4����LTX�H�s|-�ԕc^�l��ֽ:�������R&f�Y$R��NRJu[d���>�v�lfp0,c��E��
�<��#��Z&�Sz�)_�H:�:�Ai	=
�V��Zw�6Ã̏FxUu�q:5K�](6�Dq�MiJϙi1g2� J���L\VzJ��ת��PJ�uzv��֩C'V�ա)+�NF�<(���"�k�A��#�Oˏ~6�1�Y��O��^Dto��qm�r%ʤ̏����ަ��$-�ւyS�4Pi�����Q�T�6�I���9$ii��w�<˳V>�fn���z*�)*A���m�����wY��9����PN�[<CV�`�0�}�Y�Ya�/f�h��`gq�j������4��a���8@�e�i�'M�&6K �WKB���"H���,��WJ%yؔQ��D�����ȓn߻��|phy7�,FXN61lV���X�����T80�P1�#����߿�wVw�gP
Oϧ1�x�k�X�>�Cm��z̐-_XH���bc� �������>�z~*���C�I�#�ުb�=�Q�8y̕���$6�;�{У�P�pa�� U'	9��/u�5Zsa<B��l��!��QD1�3�����3l�=���!۪�*�Y�C���+̰�L�����&�2���fK���P�,���e�4ڣ�>�A�m�`�WI)�ڝZk��\j/�:V.o�����ސ�Oь%����g�Jka��&��S9bY��D� �t��YwQ��/�'�#�e"���Qny�G�(���!���n�u�ȉW*��^*��⡴�c������i����B�Fv�h�|��#�|�FGc�6Z���B+%xL%�1�b���N}��>��q,�Wo��%�e��^�^PS�Pk���n�U
{�[Y����r`ܫs`�,����ǚ�� c����I�a�ꛪ��3>K�55��>�o�UB�Us��9���Q[{��8��-NDsy�^�C�&�G�̞#SQ��7?�Y�4���(��K���Uzs��B?b\-�W�=��J@�ƶ�9��kRA_��K�f�v��Rq�q(%J} ������l߱#Oe���j��«�L'���8���c���:���gzq	٢��1C��fhSZ��`f�"�Q��<f�)���R�jP6'9��l+�M}{t�'Fڹ�uR;�/5��#q^���T�Y�K�I0����U��O��Z�������P���;����7�8�}�L�Mu�twQi����(��l�n�Z�,�R�~��|Î��� ���i�t�����m���r`�tP�ܢf����)���-vp2�f��Ss�������Z�>��ګ#A!=��Б�F9-�#�U��l�d�5`�]t8�F	�M �Ƅb�.�D��m�@~�n�]bU�Y�S��͟�$�s�`:+������Q�
f�q�0Xh]��6��#ک�ۻoo��8��r�E�͎�����<��������h�C�=I-���L���Y}�?A����x��5$�>b���[\�x~��h�B�F�AaB��J����mF��R��6d�0�"۱<���;@�����i =Ij։Ig�E���>�Et`�5��T�.lk}dT��ͦ��ɇ��8�kV(tr������C4����O-��ʋ�#O�Yc��U$��^�ry���B{M���-��������sב���
���.r�*^8W�g^y	�g/`㨉;w�b9���'�.��g��le?z�&�v��q��������5�TX�m�Q׶ R.Y٤f<ըQ��]�Y�ұ}�(豫xaȲ�Q��=���5�#Aņ항�x����_}������Q� ���<���ړ�C��F�M�zD^*#C�\�R}����̶�P�7I��}�:U2c?|bC3�
m�i�{s�קTF�G�W�J��A�7�Tt�H�<q&����1�fAXo3��">Mx����!^����Ϻ�D�S���>q4h�a���#<�Fh's��e��dH����f՞�#�Hb��`���f��~��rk[&;3T*sȱo,LMc�푫=D����md(��#��Qa��	d5�I�T�`�j�KY\Fo�FT���y�r�/�;��l�.�;(�6��,j@�k<�����V�T�d����}4�)�e¿�$���)r|X ��xFќ�S��L�R)����q_[kL_���-����i�SN%78�h�[�9�)�`��&�y���7`i�@KLM1MU\yk�L�o*W�|)b��$�(�I'>�J��%�b�ABz�C�4�j����a�WE~���l�=�;��4zF#*��Ùi��Y$km�_@��ff���KS�9O��e�N�1�P�츃郇(��Q9��|}�&+�M��A���C�CJT��O��:W�R�yqLϊ���3k����!��o~1J��9@J�F��{s�� Â}mz�9����J��գ�`j�;���C���HnPں���M�{(�'#����u2m%�~֐1Ȑ1%����\����ַм�c�n����7Qؿ�Rk%}ɛ���u�2ƹ2F,�����u;��I6�HQ��?�d����I��Y�#J�"K�0Cܹu�.�	�7XL� ��$��@B��4�}�4��b�VJ�!M�����E��Nl3�GȰ�a�؁���UZR�����x����e��f��R�Ҏ�˱���ɲPpRX�m`n��1{�OP\�������.��H�=�"���)?{hS���Q)-����h0׎��js�f'�Y�1��~���0��h�M$6�@f�C��6P5���,�F� R�Jd���8�<��@��v(#;�E}D�N����6J�U,%�XI!Z�{{[������6%
r����l�6tݸ������6F-��4��~����n!Q�¸�O叴������;7��qs�F�i��һu�6�������>�=�0�v:X�����y���>ڛ�l�-l�Q�[������f��cI�!E~5�W��6�p��)�R|y-��uR��>�CE��T�i
��;Eeiz�-$o}�K�x�]��o"�{��ҲkF�!��P��3�)Ґ}��`��y�M�T�nb��.J�?A��70���;2�\�!**�	
�N���)��ҷ�(���SlӠ����������n��>[�P�� �Q�è#=4 ��H��sJJ�6�ak_D�e,�9Q�?���e���lV���	a�,�@<���)',���'�ܬ-CKO�E�7���"E$ʱ��&��� 0���}�d\>=���c��&��H��p�C$v�C���̶�N,�)��0��A��s�Ga��;�a.�b~���!*ko!u����C�{�=���B��R-*"��D�V2�7΂��,��h�����ډU�?:�F<G�6����_�I�/i��E�X�
�終��k�@��������	i�?�"P�Ґ�mSѧ�D�d��T��~�JP��<���f�ڔI����p}&�e��c�=<��E��҇�TlR�Oz�g�L�@�ij͔�bUK,[&=�Jyb;�؆�7�=�7���`p��H�~�Th�${��cq�1���+̳(9*�;H���g3H�(���"������;$��&��|�{���'�W���(t1�"I�h�����G|:h��^Z,b��<X/��Ƴ��"����C��I�9}��e�/\��IA֛��[�x�́�QR����rt��6���}��m4���V�IS;O�k�������Ρ�g4�Ł�̆��l��觥��y3�#��&��nq��E�h��>:�}y.��L�-�K��i�]$������9�.YhZ��G���Q�aV֝LVH�5��T�`q���5J���:h��0UWQ�p`qyOab
���Q��U�,#��Y�G��][��:j7�I��	Π��I{�U١�����m�c�/�CB��;{�G�،�����kՐf��w����T~� �u�[Gk�F_��ۻ�J��|!�����"ôl!�x@�J���\{%�Y*c��h��E��N�~�~�J5�.�0E�,[�&ɴ�B�/��������#>�)`;�G�Gm��*q-L��88���wp��=�>|�*�f��خ�^�����V��� u��D�8�2����{�0�jUZ���
���>�}�o�')�z
�&Z�:�����7���#�i�{�C%�����u�JW�
Z���?6v6q���,{,_�
g�4C���/�=zPۈ���V�jt�٠D6�P��/9l���@>���NY��������-tk;�v��Q����c�)y%_9���OK��6��iZ�ZoA�5����c
��Q߸���TkG��Oz�;a�U���Η(���2�S�D����۱11"��U�A��ӷǪm��C�ZdO�.˱L�U��>h�o����0�)h/'�}&�����n�^	���-�G�U{�=m W��?h��͐�Yƀ��W�Q�k����㐃��A�/�d���md;8���`���y��s�n}-g_J�6��6� ��������l���,���Wʷ1�n��s����ڝ�E���4z�*��[}{�-�u���؆9��mj���E�Fͨ��"��#��,�����4�1-�orW�W�A����J7��n�q��5{�RP	�[��!�h�R1�DRk��&�9͎�1�XhF)[*Q9LbP�٬�H
�ޚ��o�ʘ�}6H&�l���F2N�8/)c�D�5�Ÿ�GZ3�R�(��3��0����~�?�z�Ǥ�쓽z�Z��.�4H*40��"Z�i��S40��62����}2��lb�}�����}ջ�A��<@�cA�JӘcg�F՜��`ԧp����^���}ʬ�7_\.�|)<��{�N�w�7��G�k�\�!>���P�
����Q��?������C�h�_.�p-����h�y����H��K�1D��@w��d�1Vfx�/��.��fä��=�ތ�q@LR+/�J/��	��~���}��͓ѳ�S��x��@ӦM��dl�3�^�A�1��������0$k�<iG�!��2Q'_����C}�s�/���4q
i?
� �%�	P�� �W<�Ea>N�24?ݞ���8+���<�n���;k�A�v����q���B�;i��c}���4������jXn`��.
��c���,'�B���]}��z�f�z
Z^Z��Y�T�S���,Y�>%F:Q� ~��?Bk{�F����^����v�S��X�r�o�4˫�AD�eIh��֓�W�c*��qa��z��w�t?;7��jk���;x@�vx�^G��$�iQ�������&�ɛZ�)��I������=
Z� ��Ty���{Y�����q�F��qpD��i"ǲ�5�O�i�:T�8(5ZT�E��7��P�6(|G,[�4+�/"1w���ё���C ��U��y%!��>��s�����N�:;la�����6�7��}�t��:m��DTd�s�5�_z�(R�I�V�<��TO��:�d*�H��}�h$}�&���/�g�Fҥ<R��mSPm����C��X/K%*G�8�ш�Ikz����	*����V�}���g9h�7����TB�6�Uk-A���%�&�h4d������b����$0�)o����I|���dn<����`����,�}K�/�1��i�Ioq�E2:�Bmg}@R�I�h���W�:�a�i!�������T��1��Fu�>�5*�#}pv���V�v�V�4�43�aa�9R9h����̗G�ti���]��=������Rg�>Q;���d\�2c��
z�)�oɪA�~���엚�	�A<��R|�J�~�Y�Z�Rvx(��/�]�(!~7��A��c�/6>� �y�{���g�Otg09+�c}Md�D�`k�F*-f�-}Ic���(?����2mY@i+�V�
����SP#�=Rz�=Tβ�]B�Q����ݠ���k�ӎ\C��//����N���:M'�=��1e��l��i�,�)��Y�>��&��?�k7p�O����M>� ��G9�Fe�����f�:?s����)��M�{���B�,�p�D�e�>$�Ŕ�����p*�#��6��D���w|�Z���~x���5�F{���^�Qs~�!Vﯢ�� SZ�H>��Wmb�Q(&.Q=��ޠ��+�1�O���{TzRy
n�6�~3��(�~�֝wi��QO��^�E�u�,�q��5�uP=�5�CZ��G�͜ŀZ�>b����|v�����?K��C��AB�� �> A*,�ib�:~�I<�Io��.Խ��,���;�kLŒ{Ą:�t��(�g�!U�ی�����
r��UX��/
'��[L:�
n�ɮC�6>Kzk���Ǝ����Z��6�) �븐��W϶���B{u����c{V�th�h�?
��v�ixM�wt��<K�|���C�-�1jr�B�q	*ĵ�[���Q�bgN����왋�ȖT�
��T�4K����ϢG%J3�>�$�"�����1<M��;Z��Řm=Ƕ��Kgq})��[�p�V5�H<��i}i�C�r�B�>�¶�K�}����Jj�L�I�\.(���鳚Nϒש4d��KZx}�]��k]Z��i�g{S����D$��O�^o�i�ħ^~/��y��"����z{T
�-Tգh�8��Z����BVn�i�%�Q�a�$���q=���VRȍ����M뵂�)�i��rpN=�2�J�k��_JY��'�7�M��#��������xw��&����PYXZ�է�Fen�ug{R)�<�F�J�jy�)��B�i��5y�r���Z��+��7V�H9��ɗz����h�=Ӳ7����mh}����P�?ZG�9���OnD��8҇s|/z�%�D|����?�� v�]?Q����4۞�V���tg��U��6�>]���;l��+{�5$��sT�8��V�#Q�dvT��d_
v���-�ru
/\?�^��[l'�C�vW�V��Ed
ϲ]/�=9X?D&W#����%���O9��B��q�&v^�Tw�JT��ϙl�ss�z�)dX^�5�1�o��_��,F�KT��O$?����/��� ��֦��G��}h���3/��]Z����D�I�&�R�)�Gmd��lԗ�#��tЛiZו��h�ȧ$�)۪�Π|R?ϐ73���BڔY��Q��A@��o�ѸW��1�7���Eʅ1�AB��5ʷLu�b��K5,�dls���}��1J��ѩ����R���2ΡA�W�c�e�P)�eg�+M!K:d��b��������`�ƏM��9�f
EtƔUg�>�R�g�}
����"Ә_��`
M���{n1�O-gpa*�E�?�V�.A�n�?}D~�b��"��J>�،E���8--xK����P�mc���J�JPy�وyY�ra����W���
�����{���L	h�Af����$6(t灅�d�H�
���*���l�ȧ
�T���� �����9��
�@��.��K�ʺH�JN�)p(�
VQ�2L�Ud��N����D͞s��L���֝�!�H`Ry�#��2a�4t�t�JqӉ9���q�(��.s��H>+l|6e(.�����u1P��АJ�v�����J=�Ԭ�^�Ub�ӫ���<���mВ�`%ρ��T�˒P�q0�KYТL���@;��-�_A�����G�H��󕂛����TriY���W��]���c�xH�IQ��i�M�#���mk�T}���@����5�2��9��+ҦH��W�Ԇ�E��U.=��P�l�6��+�Z4?���C��噿�����5���_L9*��X,-�$��RJ��*Ӷ�����LI�yLOOann�R��!/�,��Ҋ̚�Qy1>Qv�/�����8�yc�V]IC* i�1����p������q��4�i�o}= 
��!Pߡ�6� @�$��2*��(��։]�G:}���u�K����k�����h���H�,7�L���=I��-�|a���b�?�=*�>��Ә����I�\Y�E֩�W[G��KE�}���Q1ӡ��7�^C�o@�9���J䱢=��nm��~�#��~�-ì��ʯ�$�A��g��(�ã�@}]BR�I^�ůǮP�{n#��A�p�\E����f=E
��R)Ki���v��h��3���)>�5Y|�K��o��7p�闑%��J���C*���<����s���/1����*��m*o$�Th3�#*L��u���MّeyX0����wyi��Z4ޞ��G>��͕�d:u뇐�GW4��ul2>�T�de8�f���o�Wx��ѽ��]Fq�����Ǔ[����	yۣU��먜,�� ������L�C[�P�-M�fG�>�@�N��e|�o�>��i�f��nN?۞�f���o6�c�i���K�9��,U!*j���deP��6R,R.~���%$:46j���oYo�j�A��-U����{���L����Q��1�X|�7�;�[�u��Y��3�R��4y0���h��3e�F+�(���D�Ӈ�8Ǉ��/H�7����d����U��ЀmC�����o����ڎ�}r��!�x�%:y,R���-�����X����]�M
e2CK�o[�P���q�
�B���`q�a5v�m
S}�:�}��syj�̳�u�]E��+�L��]��sʴ�z+�J���H�iYe�����6�I�O57�m�	;�1���A`K�ڢ���$Ĝ�3B����&�y~�xQ."�����nu$Տ�-�����z�t�2Ɂ�������w�Ke�ը٣�ǀ�R�(Y*h���w�i��Sx{h�1=};.�^O��jF{���%�x�n�F%��QkP6(�ͺ)�*�P���h�{Ԧ`?|�t}i�f�/��7_�x�aM�x��d+�>���,>H�ST	t���1��?$�J��7ۦ��,Y���>��f�$ܵ�H��"!�+K�L3P��R�a=ӕ��<KaW�@�����q�#=�d����1�<f�5'��ڂ�PǥD�ۋ�;}wR�;��f���6��;���݇�Q�u�hw��* ���4�d��z��iQ��d�Z��e��=���uHŀ���x�G!��5�l6p���&�r��E��7�T����M��۴�k����"�[��5������.�C�
l��h�,��}V�{)�)[{G�����(4�l,1	�'�ա�t�)I�a�y֯B~�*�o��!	H�a�lk=C&ϧ�-�ַ�:�'O��IAn�}���Tn���k�5:׵[�/�=����d�L���`��ʹ&{sL��>D�c�Ò�%#ҿw��a�<D~a��Fگn��hq���ݵ��5ەe;�0.e8�w��mƭr�F����-Yfj3��V�,n1�x^tyr�.F26�5�<ŏt�>�>��#�􄼞U�
���f��b����p~�mD�-=�4��h�4c�4Z�P��QUO�ۉ�����7T��lA[��=�]�ZG-���!�}��Wٯ�Hi���3y�d����W��+������$:���Hsfڣ\c[�l��׍O��*��RrGl�=�7���v���mv8�Rv�)�^�cv�O�k�MSŢg8b9v�)Ǳ���<�ӕ�<�#��L�<�������c〖&���֍a�!���N��j����ڴ: �H��u�u��������c,>�,���������ޡ�Yŀh������RK>B�JZ��@��Ӧ0i�j2����(�^Co'i1-��v��S̒y��S�����q��
��hy��^K����+I�!�}�$!4P�x/a�AS�,]H�����N��W7r�}�(L��8ѯ��#�8��[�8�S��Q�7��-���6��=2(R���l˥z2�=6��I�i6�}��������M�����U'��|���D�D%��ܽ�dw����J�~?�BłV��~�BV��֪T����o�
�6wyT�nw�<w�`�jV������KK���B�����(=�n��7���څ�wH����=./Oۛao�D���}�W�KER3>��Hb��jk#�h�{\���r���5$o���aQ�Q���d�ɗ��!�]"�N_J�e\E�G�1e�Z�R):O?}���po��}m��<�~��f ��Pű<5ͮ*X�٦Z�*��W�Yt=�7���v�bkm�m*9�F͎őn���Bfp��-/k쳤��~~��	C�y�[��Ÿ~��>�u��T��l�.�|����~J��e{�z%��\�V�����I�kƒ��o��.��K3J���տP�p��L��-�^n�6˟������̑Uu��)� f�%4'o�{��џ��SP�ɵpq� �{����61��ِ�INE�{j�Avv�T\Z#�/�0,h� y��@V�2(}BA�p�Fw�ПYĀ�l����}?���`u����0��~Ѣ24�����M��Zo�8����0WHo���yt��%��&��ꬽ��7įu�}�Im@�ў^�y!O~� [�1�OW���o�Q��~�R)�����~f�c~�.F'���IW!��+���ŵ�:��ԟu�_�e�8<oT�R�<L�b��f�/+H�AF���q=nMu���V, Ӥ�ac�T�RT�Ѧ|=d��l�}��JM�n���g�1.�7!�%D���e�!�%)����ؼ{w�cgo��O�7�)��9F��v�	����܄>��V[���M��r���}����y�����}���K�c@����ڷG#t�|X��}tp���j4�6���T���1��3�xqe
*T�H#kVQQ4$����fMq3���H�"3���T4������ �|P�v������_)�@��F!ף0�E2��S�SH�[��d�m��q��P��*�T�z��0nԯ��5W�?��5*H���4�)|8xRf�J��� �M�pn�"�W@��D���A��!���v�˴ �УӀ�`:G�2T44���C����25�:�J'(F��"�p-g!�BX��#$Dab�4�_t��l��uHCa�[�S�&�2Z��U;z'i%��ѥD1�X�`Fo�Q@P��/�z�h�'5�@�1`ەs	T��&-Z_l?�$L�8��62�Ud:����
���Ю\A;�H!%i�A�B�ؠŴG�^}��;du�C"e��9`Y�Sv�m��0�/|�+���Sx����/WA*[�v�:K��#�g�,�A�h�������A9աu��^�a�Di]i��:}[���HfAZ{˂�3��7��3�c2���R�kۧ���OJ�YwP�#H�2^��l�>���]{��)���O]E~�n��uXW1�A���2�JqY~��%�c��9 h�g��dJ�C���E�K�u�Gce��&���I��q�"��1-X�e6E�H߾+\Bo��EVD'�&E�f�5>wQۼ�f���f�L�b���>؞P*�e��x��}��`yn�:T�hB��&,����<�������X�f�F���
�ZSB��L�lZ|O���jS1�A4��&v�.�
�C��C�(K6�����
!����Ƌܞ��zDE�˘.N۷*Z+E�25OeP���6RGGHӘӣ�Q�|?����y*ZszRK��Lc;�>����������~H��>6��.Tl�r�]�O���L�W>G��i�uxx�qK�ޢ�`��)I>Ҿ\Y�B=����Wɍ��gi'�(���b]�y�J1�g��ע/��M 1q����K����'�鞷�oa?�|��L	ӡks�HN}IN�ci�RBH�$np��Y�<���R�i6[�5=�1�O�J�Q(Q�ࡏ�����<*GZ�F#"GY��f�	��
�ײ�1��T��Em���lb92Z�Ю�4��M�A�{��+�}dy�c�)�0�i�TY��-�GfF�P%���D��五���]t��0.��0��P�R�ޘ���/��_����!J�e����y�t�J��I���C:�D_F��W4����	4>��1N_Q�'��WU���	����Ӧv9��I�`8��׾�u|�k����t�=��D�\��
$}b@�).�3>��Z=S�����T1���,�
q�0� �}~(2�(I�K4���<�1��4����[@(�Q�R3/R81�<�}���UJ�[�0!ck�r�d)�ӻ5֑��^}eؘ#⃍�A6X.�4�����<[�Ƶ�3���	����O~u�DqT~ݙ#Ϫ8({�H�?��;7�/`���`��5�s��&���ձ�)��U�S�s�hSe�İM��zC
��^Ig���m
��y$8�2}��f�����$�L��rFBW�R��&Ϊ�!h��2MY�F),,;���~�F��.����["܇A<(8q���4-*O��d��C�z�����U�=��#<=���l��
,å�C���xX|6�)���	���bcm��T�Q��'領��T��[�,@�e<�3�ԅ�0��6�:CE�"r��P$Ӛ1���2k�C�[R�sC�K
��d���Rބc�,�X=%qi��STƵ�8I%r�2I֨��1��.��<�<V�p��5M+L������b.Z[=B�j�ZD�N2M~��-c��Y���HU[(0V�L�JIbc)=��n���̙^|L�����]��Gq,�x|"�;9bX����<lSB�A�f�5k��&��%J%��Ir0�ME��&����*R{ZzPGB�,�P��A�\F����wre���m	��2e���<�����1�����9�R��$�f$����TlK�Q^-f��PJO��
E��B9K�<ƺ�ȋ2�+sS8�<
�it)S��JK�C�f�3B�2%��^X�OO�@��i��j�1̕՚U��d�rT�>�ou��|�.�[�OC�
'O�Ӎ:���v�6�գ1�J2n@Y�o�Yb�.!2�Y�yS%kTL�?�E$��\�a�lC�}I١E�lE�,ǔԞyhIC�
e��2FKWљ9��t)O�74�DW}�����vF��R��5{Ȣ�ko�j���
ӈ�o�2���e�����͢��cz����f��K��Y|��_�+_�<��%�S9��4�4�(�H�iņ-t0_�RᏲB�	ƭI����!����rPZ�����u&�*`\+�
���b� ���=|{����4W2Q��/>���y�=�s�֩��zY7��Qv8MU�rV�F��<G������3{Z�]�Q@SKP���&�+G�� ��*�-��xCZG�Y2Hqn�>U��2�g_�p�)rz����83�X��-E�A��%�8�y6	��8�di�ֻfv\�C��,&ur[�m4 ��Ǝ�$ᡛX ����!l�n|�k�ti���x���X�Ұ�4?[P��X
��F"R��飷L����$�*����H�>7͠��}�NY�R쌤��2
�r�����Қ	=Bc����Y�Q��a�*�sgК����S�%��+�zр��Z����n1A�,�$�b��JY��拾�Y�)�X��}-�Z~ə�LN��q�(H��a��{Z�	[�2�NxK�!���b6����7P��.��ڋ�Z'��^�7z�Y���:Ϫ��>��HQ�*�J#m� 
j����y-I�R�tH���8������_~L>��O
L��p�7�.���~���>f<���{R<钦�.1-��)	lZ�Z��}i� �fj���Bs�ꛫ�w)S��K���)*���YWm\
���Ef9��\�0���̛��d�m$��lǰL����1#��)�mv����{�
�,֫��Zy����)(��L�R�H՘��`��Тo�0�2���i�nz}*M�)}z�e��G��P�B�� P[�F,���ښ]�#Q�lpWó�֋�F"ؽA4/���(-��Bl�B����*���a|%�4m�����B�m1��
P������7h�Z�
�k��@��kPrp�_>�!�I��̋uч��x�D{�<�����Ic�N�K�@��F�Zӣ�^>!-�h��t���?��9S�4#�ͮG/����w�����,6���`43����^x��,,`s���.i��	��.�?(_%�[z:�<D�I4b[�#�������g���aaM�����.<�,s��Nv��0�Ҡ����E	?�ѥ��02�K&e��q#I�ϖ{P���^y�N����խc��Ȓ�i�$C#�v'O����@�},{���"�Gv��d!���6:�C����If��S.s,��{*ܒ�,�G*bKϢ7�4R��1���<��g��1�f����/�/AlmAyU���x�W��e|�׿��Vol�P-\�2�2��%�õ�I��R���Gƚ���Uq�Q��?��jR�5��k�{V�6C���M�ӄZ��Ǽ,7			# �6�#���.v[2�ܵ�b��F/a�ֻ���{��(9h��<J�^)��Y2��O�?�j�ϢM���e��h�p�Ӏ��r�~����6�lh� o��C���)<3�s$x�Bz����.ct�evf	}�t�g�iQ��I����B̴�����Ȅ�v�fh%䣁u�t�B-�1��:�:���R�$h-��j/$�d�I[4)+#���~$.�Pb6m,w;XD;+�0��?ؤ�>VC��N"���qé�RHX�DH5�跪�cZ��Jt9�1\J��%�y�5��lK�צ �#���֘F��/�L{�dhͦSyp9ZP�|�s/�I��ЦmRp4k�]3I���@r���w챝� %H
��()�y*���1��V��E$V��r'!-eM#��5X�4)��?�ٸ�F���s��D=���qxxhk��٨����btY~j/F�����LyE|ځ-� �� ��.�<�]&<򓀵�e����!m�����J�G��
�G��6e�g�a8���r�Y%gp��S���#Y�Z�:Lا��}���)�i��ۄ}��s���ψG�Jl7G���Β6��҂V5��}{R+���JtL�
�?��٧8�_ư|�I�3"�LȐJ����=����� ޣжO&qD���>�tH�
뒚]����}�w�i��0?Z��ǔj�Q����-�ת�� �_G�GfCߋ�EV�/�K� ��0;��+c��g8�����@eN<�OY��47ꪶ�M�f<v��]�6;��IH��Y[���mA���/Y@+^���x8X�8���䩀�[^-�H�Gؘ<9�bcʟa��W^@R`��6����tYO�%)IX�|�zk�JC�`�
4�V;��x�:Pɖ� *\��+�y�
�33˶ﲬ�z�g�7 �QD���B��ѥ�3�T)����r�������A�|���eyfɛl����"�S8}�Z�<��aWF/�i����R�!8)m}��A���C�<�q�:��<�{:<�Զ��-I��뾇�p<��1X����6�eu�Q��T���j"���4�R&�2���W2�SG(K( 4��e[���"%*8�K�M*R��ՌwYOe��{ڨ�+��Q�x��/c0�4��瑧1�o��)c���)ʊ~��5��42�3,%5��?�����=|��>�F��������ų�@�r�2I�X��e�D�q�Rc��Oh����U������q�y�:$�h��#H�T����ݳb6��ƈ�c�Jrg�����%����7��c-[f*6�aE�4iT��cB���9��/�E��"�5��a����i&FhW*kj�2�i�E[��>1����4z�gѥ�<Z�L+w�� RL�5N6��{68���fA(hF6�32���ha��5��bW}HYo�hߐ�����[0)ҡ��V�������R����_�R�ײ�n_����Łf�u�!7�fX���m��>�ϝ$�钴dSz<�:���ހ�y@+^u��UZ�^?fXW�u�Zb��N#���[�TK�B�6����U��e$�3�'�O�eE���+i#�R�[��H��1�Z�@��>�Uaq-=����{�<g�d�ـ#��BLFa<�9���or��ͭ`t�2�Z��:i����:����!>ce�^��ðR�BۧsOzIa�c���%�ϑ�X��Qg�5�Q�E�:r�A�;A7T�z��c�����@I�B�7�:��m�{�$F��|͏m�8Z`�Y��ȁ�-��a4{��6Gi��F-�Q��-��x����0����1H3����ަd��l��
R(x���=e8��F�ᵿO�m���3�SK�l�����$�H�e�E�~�4���U$ο�4�4�S�������ӬȀ��&�{;UAs�
��%��mGZ���i�����9ذ�X�|��_������,��Н-����
�R���퓯��\��`yɫҳm��R`=�Q+d��y�'�� r?��E8����~)�ZH�<��Q�xc�嬚,�e:����|�g;��fz+�@eH�����@�Zm�3��//b��4RW>���UI3l�$r}�a�e���t��m}*ã*=����r�f(�h��^V�E�m��Z8���x^��s�]-S�`�9�u�������
*y��g��ǭ�H9b�d<E�����imc��Ĕկ����N%r�m�{�s��!���r��#�馗p�kX���Ԏ�E2��GMt�TG�ʜ��)��\�Z�	�^1�hd.>Ŷ|�sWh�m���٦��4[� @�P@ZK\�.Q!�F�c�o�z���T��Q����4\��Fq�2�T�m����ϝ�S�T'����UܬS6�P���U����īh`��&"��<�&t&_F�S}�L�{8,��k�q�c���H��f���ǂF�yH7A���������=<���#pPF2�]���ء��c�9��ÆNM�����-\��Obp����_&g�z�T���P��p��(�P�`��D��RZ<�0Mm:�E�	ZPEZ�+0x�S��_.~����C͐�%YNM+k�CY���G�`�i$v7���>r�LO�m��-��R=Z�md��P>�Fyw��U�OE�;��8ZR)�4���<�`)�r��v�m�\ʓd
{�O�t�%nSL:ķ�W8��ő����]�}����Q�Ѯ8�A���ھ��*��&d���j��R��ZE�p�̯ا�s�G&gZ�j*fc)���#ӧ5O�-���5��4��p��cX*F<2lO�֠�6.҂��۽�it���=���nP�K�D���$�rL�= ��������,#���<Z���2=UAv��T�ZW>���W�瀏�6y�?Ͷ�i9�H1V'g=La�"eĔ)$�1ί�b:�Ý�����.����}�^��z8�r����Ukp�m�P�=ÖAx�,��p�)�R�F�;���]��aA-��7�F)w��2���*���L�a����a���~�6��+�#��Ie���G��D��|ZE�ְu5i���@J�r�;�|���A�K�,�q�N��0�����"��א?���g�K,qP���@~*��;{��]Sb٧��H�.�����ʖ�g��������&}VfV�/�a��E�l�� � iFR���
�qFA�M�C6�E�*M�77����8����ǹy��Fbg5���ۭ��Z����/�O4˸QN��s�E����.>O�*�='r��i�;u��
B�[�<'q��� �[��I��#�z:�}�5�vX��z�H�|�W[eLJ'��1�ߐ�@��m��\/
��<�����䖇ݟ>;�$��v�[�F��^v���ZR=�q��C�������&b��sh���;øy���Tsa:|�&�ZP]�"�k^!9!� w����ߵ|Nfʡ��]e���"}�j'V@�:zk�`p�Կ�����C�c*τ2K��������$��@��t���L��A8�So��E)���+���`A��W���)��͙)+1��]"��6���d������6;��[TnY�r����Yk{��6�C��G^�O���0���k�`� ����g�H����;���*e�m�9�W��)��b95�{�4;V���̰\�4�c���Q��f�F����Iʎ?�h,G��sJ�`��er��Σ%ҟaFԟ=����/T�,G�/>�� L��Q't�I?mlz����_����c셨w�'�(����x��Ŝ7s�&�_&���h�6g���C���{~NC^�������ͮ�D�z[���o
��տ禦'˾4���8:�>!���?Uc�v����g۸���� ��T[4�$t��"P{ _s��5�>����Ff���Г
L���TD��T����N���T��2�"�����6�j�R5s�q�i�/���H �~#��ԇJʓ2L镭U��C��U���:
�a�ts3A<���Ѫ��λ��Y����v�'X��_G���������
��_�
�����H#��4�U�Za����)f�}���.�]���k�7U
ģ�iR���ULͰ�/�q	���7��>��)^�v1z?��>>=��Q�8ѫ������~����~�F����oc��AC3�a���@8�!�z����.�(3�QՊ��1*=¸��rSM�������q���fCu�H�V3�6���F�Xj&��%៴�������p>�u �'`��({N|�eF���Y�U�Czn���e�ٜI�i 5�ǼPAzud�C|����[����k�m� ����=ơN�W�_A�����47��x�~�.0��4<,$�cR�X�p^�Lu���*o�W�y��!ù5�.��Ģ`�LF��T���`�`�pS�3�M��o<0 �8:j�S3�����Ss�q�B"#��t8>�-�rHC�lL�i���Ǥ���D�T'��A0�h����N����|'��/�
���Z��I�0Y�a�S���F�G�)=�bo#��"�Y ��h���!ߍ�L[�G�KZ��tJ���z4�!�:d���0�2�=9lB�2A�����1z��Ͷ����G�����]TF(�[�K���#������1����Z��iS��O���<���#+8�\�g}�o���{�3�H��Y�jD��X(�K�����j���w�v�N&�z���7��M��d���}|�SB����~�$ �(��SM�9R�Q}�嬮5���{��#ҥ��Dk9��Vm�_ (ڠ34
|�k�q��F{4b��x�y����>���cx��t��� �(��n!N�����7�A-#�$��M5궉�BN����'*���S<��������D_{�����k`�޽�n��K%{�57��'��4���n������J������(����B� /GF��6g��޻�{{���#E���q�_|���q����8[	�E:��Z5ãf�頧q��
����`9j*�Q�@� zH�>P����zʧQ�"8A�P}^��	x�O�<O��8Ե���)�]�;B"�%��6I�N ,�,�}ĲV-�㗬;��r|)�o��І22�mtcX�JW��u=&�;1��J�<������v�d�����_���&����R�q���*�-�����;-��i<$9�NG�/6���hJS��(��M�O�:m6����j[(d#*�1A�G�f�A2Z�F�^*)U,�9��j�ҳpf7��y��Ĉ��	"z~�H��72��#Շ�G/T�0��6�||������Ϯ�g/"�4*%GXHy�4���7��U<�A&�m�T�9A�����A�v
�@C���G�Fip��9��Z��3���5/]s�����u����s�A����w��������\ ?xa�~������C�教f�C,ƀWn\�����}�AM�J�tB/�%���G��Q�j�H��V���a���j^�
�����Jћ�p�.!L� �a)8��
a/�#�������fJG��a�<8n'�h"o"�qN"s�3T�T
m��Ct�hEX5�u���|�U�}4@�A;w-���`腍[5$}�/��������T��èT*�&�Ѓ��j��ٱ�&k>��)��}�l�*2�4.��{62���_x�5��q\��J9�+��sNڦ�I"�-��x��Q�B���Lh�Ӫi
�\g��𨝆��	ś�K�i�w�I�,�H��jU-&S�40E	��3�i.J~��Fx��R�+�fPV�5=HFi��z�24�W�dD����8��h�GfW0Y�Jp��r%(�%h�� 
��L�<kZ=�e��A�!S��VQ����$�]����0�@*2��_�3W.�z����)��x�i,� ��5�b��}٣���+���b��jw�X�f�7j�܊�gR~:���ڞO�Ky��V�����b�\�K����&��SKx��^~�&VW0�7&M��������?sm�,˲Y�W�A���Rש�˔�����[c�^�{*gr�C��DR�3��6'HM"VXA0��l3\��
p�n��|)߼i�}�3y��� e�tf��J:�.a0G�+��q��y�dX��(ޚ�a�%O�C�#�I���@��7�L���ԮE�iyp3��3nr.�}{I�n��u~je�s��fɰ��Qq	$q�����{��O�W\��Mb���c\����(~��|����,��"����<�B&��.���y�{g��C�9�ыe�O����j��*�Ud�&�f�e8�R3Y:ü���d� ��@� J�TM��aR�`%������� ��G����M�L�,��CPݢ�-FS(O�L�<�Y3�������<E�!�\H��T6���F������)�"������v�q�L����m
f��e�[�V�/n�bA�4cv뜱x.гGA���.JM	4��ϴGP�,YC��<��7� _�VA���<Q��F��N��~����(T%M(KR�D���Z�Xe�L��0=��O���d4
,�ﲀ����tM�E�b ���k����UE�%&�N�~u��/��n ������3����_B��q<���^���<����(�;h4z�RA�i�'��}ߚZ<��d����s�>������}>�צE����=�θl�ר8�u���L��㕍9��/����2V�0`�*�X'px��̧ex�X_����2��x����~��1*N���MZGv*D)�����M�XT��lQh��bV�d�ZE���33|��"^������I�2��CC�r����aat�nc���K�{�o�E���(�C`5 �����d�=�&�,�	��>�}�KX�1hT����[QT*�^�`�M﭂D��5*�|���A�`T뷵��U����ѱ͵�Z�'=?�����r�`i�"���h)�0�OP�8��ܭu� �����6%+
�]ohS��j��i�O=﫯
�͜�����I��&���ߗ�e9i�~�v�w㵍N�w�\J��Y�8�"*T
��W�A� .�D���]㱅,y ����ŏ>A��'
�UQ���bc��,t�a�L�m'�����Q�f�P5L����������\�������	#��Y\ H��,��w_����ޗ��S��'���~��x��Ed<b	?n޼�|>ck�-�͢K�zT������O�iy��0:��Ĭ,�ٽ�*�ϴ?.s��k��\\�&-7�+��O������x��k�Y^E$�Do�1@�̅�X�(nc$�qĒ��bXK��%3<h;h�ZM1��������jH�K#ñf�' �#�W���\%�^$�̢�Hi��]m:5!�:���4���E�i�wrٝ��?���C���PЙ�V8�Ƃ���t��Ĩ��8O �1̝@��w.KF<�P7�H/�s�M�dX����&7��#��7��qәJˊB�Oܧ�/wsA�<���g���������z��hu�����m/a~u�EC���*��gX����9B������K��Ǉe����ˢ-���@��ō���4��ǝ:�IG�� �JW�^����h�"u�QZ$z�Ѩ�y�6���/�"[=�u_�}{�w�k�Rg�	�����n�&o1�fQS�K/�.���n�H��)DF�7r�N"��i���g���S'��ùWӲs�\��D�����������qt4��{j�PM�A{��گ㔞��Q��XX�#�Q�ҫ����|������C���Yo�r���A��V�b��<�yY�͏���c<�=��:��nƱ��"�u�*%��4�4�dHo$�&�ּC*� �����a�h T�QeC=gzs4�����7�O�����=9������jŲ�?���O����\a�Jp�x
�{E����rh�3� P4�G�r�m�$U[)��w�Ú�Ԥ�0�8����ۄ�ehh��\�����.�_��+����`뾵>~�	���Q+�Z,�K������kXXX���2�t���(z��D��9��&`�w%(�Ji6�� ���N�%���5���+�:~��%��w��_���W�x��2�� ޾���><)��E�N�������+������WW|X@ŭOpz�IcN�����	4_4��P�i��NM����u"��?�5QѐPH1P�7��qu}و�h�4�Bn�Y1�� ����̾�x�f��<x"]Ԝ��ў�{z�S�ո1Z�S�uTz�J����������\�����x�BOT�U��''E;��.�(�N�A{���>G�(��$IВH��1�r���?��)a8uTv��ٚ�X��O�!>:! :B��6�=d'5�h+{�"z�2��`q�p��W�ϭ��>|e6����Cx+�v��k�>�15G��iH׈ �괈�i�y%��g�J�V�������_H��+����?�A����z�'Z��t�v]��,�p�g5|r�E7�D=@î�Ij)w[(ܬ���T�绔�g
�}��끋/��0*/s������⟓>2�"~em�^[���."�0=�G{������C���v+˳X]Y���%,��p\k���.ڑEZ�<N��o�?�9��>`��ҁ�/g���bur��!��	a>�FtXB�TF�Z�u�&�걤���C�o��\k߹�Ɨ/�������3��U��� u˫K�>�R�(o�s6�CR[���o(��#,��G	�����}JO�ΓiA��.ϟۅѵ��tӵ�7�Y�����͘}�����Ҥw���R�����T�9��P��k��0�K�y�&:U<�|�;w�Q���u4��6J����a��L��ן��F�tT�p?�!D�y�F�a��E�E}"c�B����eT��.��@�v�d��:�#�v��<�B�w������L7gKX�u���~��Bcļt�t�yh���:�G	e>U�`��?�d-�S�8.�5]�Qe�Oy]��/H���g�tK���|s����D9��w�'��M���n�?�GDww��E-<���.��P�D(a���k��,�qi-����dldF.�#0jу=���j�(/��\�W	��2�z���\�x�
z��.�Q¢sF�>��^OdU�bU�6>y�J�:I�و��K�S�UZ��p�����z��Tj����~�1>����E2�u877
du0��ᡑ�$����6ކ)�)�}r��PO4��1Г��t�a��yo�{�J�vB;RI����>���	��1M5'�cl�����f����>�}�wn=�'vpt\A鬎z�
-T��}-��&6�/�5�P˧XGA��UJ�fV�N50
���+��{m������e�2�AO,�o��k��5i��up^���e�t����֬qa��4���D���*�n�f��²��IsUө���i\Mnj.�2�<�("�Q����>A��4y�Á�~�i$�dtlFw��9?3���*~�% z�Z*�;�@`�d�Zs�G�������hi��S�N��!���񛶳L5q�¹3��3(����:�w�]�&Sk�M=�Y�	����ԡ�Ӛr~%?�YO���9��a5�Ř��v'��,�H�3�I����e��dR�
 :A@�7"�S�A{�<x�����j� @�L�	�{JԄ7�7�!��Jڋo\��K7���En.FB6��c��Ƣ�M0�GPuFy�1�x�;��5 j
�o7���D�鱗��U}����3����>*ZFJ��,�:��߿�7?��;�;h�ۨ��pĢ,k���!���m�qY�,`�~����#�-�&sk)��'6]�j]�kl��}1b"�������>���;I�7��ԜbD�5�89-c���m��qT�����Jd����r�>�!��O˰L������iX�8�v�?�Jj�8Z�Vv�
��6B:�~q5�G��!P>�.# "]���Xe\X)���S���NQS���h��Pi����	�Dl`��1�6����P�)�O�Q��4����7���޳�=�O���l���YɹIW&ttO�7Ĥ�%�0��u:�;������c���{�U��]|�]�q��
��N�� y�O5Tmp0�PT-#rR��j���#�1�Yz��8�Y69���H�`���Dڷ��Z(�)�,�(�c�]x�G�u��e\�w��\Y���T�����8�#3>��H�N��1���4i����[F�</;ohLvη��a>��czi3����ۓ,��m*S�x�\�[/��/�&�n`R�^���|���?�m��%9F��Z�򵵩��P���n&�;��\{�Y<��S��gPky�RC���8��V�����M������� ������T�!8T<uz���LW��)�./�2�9ؐ`K�#�D
�1��U��ҭӀF���,�pr�>��}|��;�t��N����Z�Q4��=�v��Yy��}s����p�ѻz޹�T�34N	�
4r�B#2��ri89�`����8�r���X�NsS�[q�)�\O�&zO�����=��χ�k�c�F�䤊�	=�b����c��K��P�x�wR���NOO�𠈟����%����t~���[�*[���jU	�@�h�6R�[��3)��^D�ʃG�����mͧ-*�pp�3q�[sUh�SDˏ�\����W����*�>���I�Ʋ�Ki*mҫ�E��GG@��M����t�U�h�z�
��h�2����5�,�NFH�����������{r|�^�m�ibHM#� 3לFC#&�2xpr"xN�3�;2����PC���<��L�yOqj.*�g���i	$_����y��{3񖖔ф�=z�}Z-<;��M�`J�<���**s�g����t6�G%��,��<�	K�7�d�F�Ǐ�0<��o�N+	�j�gg���n�|�
ԇ^���������N��%��W��;/��P �#��j�NF��D<�l:���9�3�F�n��k�O�N�;+2q��7��"0?�a8�D2��%L^���w������w��{��G%?�B8��j:xpx���{�;,�����~;��4X�il3���<3c�;.����o.���V����n-�.�\���3���[xp�.���$�7���߸�[G]��)�#i�?���:n��~	?����kb?4�i��2F}S����"��e�#���-��8�?������4�%���*�.��O�K��q�H�7Kx*��~�&n\�C�Q�g�A!��L~�z)�N H�ԣբ��o��
�f��v<�DP5�th�5�mJ#�h{�>����ozʛOn��v����=�̞<���}"����w���>�uCG����v�B=��h��Gh��ثy���"n�vC�8K.a��qs�;[G�4����)^�[�Ij��1~9\j�0E�ae{B@6$�d;���I|�E�	���2Y L���u���p�YF����M\V�~u	�;_��ZU����x����	�0�N����#:��_�P�H�o�Uf'Uݹ����|2�'J�]*}v|�\:�4}|o��L�*vw�;�)7��xC����e�$��I(]���8n��@0CI1���l���#��g��D��²(F~���ˋ���?���]�&3���G������9~�7��6N��p�h�Q��o�D�����sv Ԋ�~���C\�M!�����^��8���%L��u�U't͵Ch�R�*w5��L���D�x �D��(��{�y	�&� ����nb!C؟�~y�b2�����9zr4h���s��!��H����t�$t�.��<N�D���[�XL��n����;��JH̩��Rؼ���pq�� �MCr΢�-0�L�Vگ���8E�7�yF�!���L�@#�(�a?iD��{�Ҡ�hAS�Hs�t��n��C%���*����#�����t�p� �����8$�_?Ja���B�>��~����Q�9x�7P<�b6��w���"�ho���{q�X�s�:�\s�؄�Td8~u�=h�՜#pa�՜-��Q��v�Bx�_��&'�����Oxt�=��2�5�CQ�G5F=� �����q5*}+u(א_���HEc��}a�����j��Z�I_��0�C��4j��M%ǩF�k ,�fU�3_20���&���>2�^����6�0wF�'�B�,;�"�lRI�*T͍&rH^��U�+]k�T��]�3�6ҽ3�����o. 6� ��@�!����x6�O�����u������1�/dO��'��+/|�Vo|���.��[��������	��o�b���	�|L� �ۯo��2����2]L��X#���/!���Q�˗Q���iޜ�k���E(��7F�6�%�MС$ C�E(�<�/eԘ��~�?o�Gs'H���avOt&����xߚzY��
��Ds��P0�>B�z�R4�4��j�C��H����."g$O���L"|��1L���P5��@�|��5�3;�O>�\P�����)�}���țd�p���|�>*��!��c�䰉�p	��_)�?��W���x��=d�y\�_����7����(=�B��`�
���3��UϬ/�����D�d�Д�S���G�0 ��ܬJ��?�X�T������2��d����k׵L�{�����}���[ҫ�l���5��{��?�٫���M D9k�;$��Q��.�������Ak� ��`Ա�2mbK�h!��I}��\]Ř�4o�3oQ��}�D����T����-y�?��g�̅Y��gx��q��M8��AJ�.F�:z�	>�_@+��Sa����^|�&�9���C4;B�z4�ݡcs��fz0����gf��y�4ɮ֣T���[�"�GWg��0���@t5��K�	�#��R\I!�n�?�Mϴ�ozmJz���f���%l_\M7�I`%�4dx�*�{��!��v���ē����������6��͋��@<A.KtLCѮU0�0��?��.��!ѵ���V�x��*�T�>�t4��4�2_��b2`+T������v4�+��XO�B4a��ai��M�R��Х��&
h%��N��`�Z�1���L ��4�8�'�OE���)8���֣ 2Ϛ�F�N��qWR'j�3�K�j}�+���v�����TG�>YI��p��2�z�T��j��D����j��l�4�uz)��U�,Q�)�a|��,j���-*��o���C��E@J����P�"'XP�kv�H� חB��+W	DB�7��	\�v���pZC�vwg���14JU�S���sظt��T�ZM���5N�ME��6+]4��q:й��6i��U~*NK/�)ω�0?�g�e��=�:����w��h���粈ј�N�H��R*
�}�=Uo��A\X\�����I4� L ������ �`��J5B�qvv�++G�hڢ�a^�"zg��5q'�)�.��3]7o\�l��z��>��(�J�A��g� M�rR�E#�4,\4���а�RB�5zH6	t�-�s.ī�y|��9,�	���Od0���Q�O���ꠉj��U|�5��^ p��A:��qay!�]��@6D�e��~�6�;ӪIOm*��:ѫ�ua��!��*oћi
�1�}�^kD�O���QUS�LCA7��d��i ��vfM��*�q2�	�%�-u�2�>PY[m��"]��c��ZH1�t;7��ֆө=']ya�Z�#Ъ��@��-MRYQͽ���U�{���U%���S���E�IR'�4Z5��	=�n�Ԉ_�K�te$��b5�o����k�H��Ȑ�U���,�!���.]Z���Ov�P���'�4���)��a$��ӥe�s�h{�>*4��a��Wv�R����o�B��Gau����M�ќ�'h�%ץ����eO��>����^�E�'�s���Զ'�ٓ'��twW0��V��4)������ȡ��G_�f�"AJ���RY�$5U ���
���h�\���E���P���G�
���j`�北7��r?xnK3��drH�1_E}c����A��RW��c���]��C�3��y��HR�f(gZ�==�C�K���9����6�eRs1�g�h6◲) ����|������C+�!}�_��LB�
�����	ZYYhws�NOu�ޛ��񮇟���/g��@��<0���\^�Х�G�
�Ov�S5U��HƁ1g��M<�	#�B���G�G�ԫh��1��.a}vu*�;h�EG}\�E����S�������q	x4���"�|�o��G�;Ԣ���h
���ԟ��5uH@�N%�0��5��˗��ãV�V�� �*�׃��>��ӳ�@&�9L2�(z#w�*?(Z�����	��h5�ّݝv�pϹ+O�[�Ę��]�p�����K�l�G�|��u4͂�,��`��|�$��G�1=^kK�ᡧ���n�����P���X	濄Ś�T�(���#P>�rԋo޸���U
���z����G����ݾ����%���y{�΍%�OZff�x/�S9��B�	`��D�Ň�Q���	�)�� ���E[k�e:E2�ŀ���e��^��D��5�qc1�`�[w�a���w~������N�T�&�L&��~�;��_�!Q�{�4-t�	x��?���ַ�c��s�=�!¤�W��
���#\�v��{���R*C�P�����~�7��)����Z�0]~������?�|���C��G�Scĩ�^}�%�������o`���.��4I��~w2�̘���;�->k�Q�Ы�'I�:'�ԇL������
�k���e�i`%������탃*<�GM���{M5e��� '͞�����똛�������Ժ�� i��\:�;w�'o?�)�ҁ����: h�ȝE�R�eL����B�&� �|���~�j}����U׫I�|�6���Y��4r,c��2~Ҁi��ѱ�&zH��+��6O�w�gܒa���׸�'��+��7�u�s ���KV�4t��6�B�j�C#u6��{ȯ��=�L�����p�� CyU-�t��f0��oX�2~�o�'�W��u��d����Q���������C"=�k��� ��;����r�@� j9�E�}��b���f��	��2�*�ƅu��'����b���'�Ӛ�ır�����I�!u��%�r�T���.���m�soM�%�=��3:�Q���2��m�;vߌ�{�n�C����ku:}�޲2;������񮾔�(�J�;�F��e>R�(e���8Ч��b#���w錫�]:���ax���&����/ef��|�g&�c�;E\Nz	�b���x��b��X"����+�"C���G��%��}������E����R�r�`a?��5���}�?RBidPVk- E�x|#\���l���o��O�碽h�nn���������X�o�fGm��lW8{_�� �������#@�]�����1��'
��^gMu������$tL5�18�#�)�>*�_����_�5���O��)�0�������y�vQ���S�Diܚ�n��Ұn��x�������la�[�W?��D��͒���BVaP9X6J(�����Ү�2�Tl�6BH�N�F#�h>4S�uDo���Pl&`-�0��֊��o#�fUs���oF��t��~I�{&�����`��b(�S�%T0&�3gGz���N�F[�U&
� �O�5��BN�H(�	������Zm��>���U~^��8Ĩ����x�$��0z����Hi��,�A��Ԥ�����2޽����}�ۘ������wqg�L�;��s�;����z�)�	���Ҕ��\�r��|���x���Ata	�\� OSS����Cz��2���B<j�S*1w�h�a�ƞ�tki��5�_������GXX&�e
�g[�R�~�������07��j�L�ъ�.^�?����q�&I9�a�B��"	�O������Pm�qF��ڏ�������ʫ_%�y_����
��_�
��?���
Aǘ �(�0��o��o�կ|��Kx�K/!�x�m5p\k��� �@�`R�����yć,{[�UeIZi�l��ڼ��c��3y��=�Lo���|t�^{�=��ko�o����v�c|��C����m��E	�g���)*4�w?�����&^��x2�+8=:����>>n����HW-��C�|f��'d5PA��2���
TK���_���	I0��F��dz|]~-a�5�ԏ*3C�0�tJ.�FCMJ̼C'��s$�ܬVW���q��ୃ
��$l���4��#�|�h1�=1]�s�{��R'��A�	÷�5�{�ޙh1[�uʞ���[�aS���0
 ���s���z��!%�2P!oMy��֚��b��M̄�7�ڻ��/��c��Y��ů�r�V.8ݯ�ݭN�yhM�q��Ç���;gM|�s���O�����+��w��[�G�V����+����l�Q!o��=A���K9W�%V�#��S�y��<i�0z�{
(:j�}�[�w�YP�ނ1^�=tO�,�1^�)��܂�a��u~mq�J�Wi��y�]+K�������nҩ �*ق�ʤ�����h�ҀF��0�����%7�N���S(�k��]L(]G:�zC4�gm"�-�tw�7o�o���ϊt&�Jgt-5C��/vk����l��"�2j��?��>�����[�X̄�h��{X��?����&�q�F� ?u��CN�-K&`ȴ]��A�Z�rFz���Tn���|3�=�$C��g���O�;��y���}��
�tSWR��+DI3D������]�d�� ��|HE�����l���Gx���m��z]}S��t��*��.>f|��
<���2��pR)�F漣��Oj�Mps-�������B���[��<��B�(���Kt�ˆ�R�Lg�`*_p����ќR6#���>�c�j��Py0�Xc�Y�IM"��[ˤ�u��Wh���1$5����	�S��8��PL�-��i�:�=5Ґ�T��!��T��kk����`��(<
'�3�20�t0" ��W�S5�J���y�;�����.�������'���὏p����w���Ao���A�_��S��x�8���[��jc���G��Y���˗P�r�������3_q$����4��#�2�&���qT*��?ĕ�jv���?a�h�����񕧯�K�?�0A]��A� N}��"r�0��կ!����L􈩹���ق�!��Q}[~�K����܂-l\b����g&�ͧ�"�b���a �8�Q�[�\6�K��T��T���M�w�cuu�TK{]~q����s�7K�䵝J��֐0�.B1�y���[&���˨F����(�������`'�c4j�ѳcWQ/�"3�b=�Z�>=�`�C���Dp����G�7*�w�p�>���/��!M����.��l��_f��U�T8N�O�K��j��<C5j�e�Z�~^��$ H$�(��0ih9D�傖���"<Q�8�a�d\�@Qnt� ^�0�6���D��ҟYc����sA�d���K�XL�tnJ��v�ʱd־`rK�C�%z#�U.C�ٗ��_��C��ahU��� A��v�ӑ9@��#��ҷm�K�G�I�)-����`k4���=t�'(��9<��K��0ŷn�Y���U��PMl�<r67^���V�����4qvvb��.-,�I`��?~�n7�/��a����zXn�Դ9ʹ��͹dTri1���Z����]9�(�G�r�sUi�����}�� �TW��οi�J�O7{6=�9��&A�������w]�!�ykD�G�$�N4�_���K�䋲<Y��^:��(�iĖ�rR�
��x�W^��A�[�(�N^�1�����<��(J����!*��{g��H�_O�!���~~�G;�Dٌ��w��=x{�������z��5�Aۃ�?�¿��[L��"�@jj]��i�D������V�����0��n�n��������\��G�Xܼ%⩨�P%��	~��B��%�1�P𭺓��4��4Z�����/2�iV0<�é:���v��c"b'?G�N�K�s�����@�����Ng��x���=����ddRp�?���jU�dR�Է���i���&/����4ǔ	e���N���ć����	��)�A��i<
���o���?ъ� �*En��D�uJe�7����zߎ|Q7e#�{�Vz���� ��G!e�g���X�R�Q���HGJ#A��>�)Zm��we���F�9چ���W��V��cO�X�YyR����#��>	g&K 0Fy��q�����n�
�t/˨������	���e�KT&9��:(���Ҡ�{�7߼��7�"23x����?��"Aa(G��5z4u��-Z���|��z�O�N�� �4�u�{ŝx-M�� 8l��}@�w���\B��ԛ�x�����!y�K@���B�x
o��1�~�]엪4��M�� �J�z�7?���qe~�ۨ��agg����P��Ci]��f���჏��dF�����>��;8�>Ň>������N���{���x� ��}r��#��}����	����^�˫�`�!�
y��]5'6Y(��-��]�@͝2䏛o	��kOR��`K������G�c��p��&(l\B1<�׏�8�Y��r9�h�k�6z,�VĀ�7E_���ɧ��7�Q�:�����gIGF2����^��) Z�bB��N�"�f�tܦ:�Q�x#x�]�����:4`��(Iv%`*�)/����_ %@P�#����c=���6���d�t������;�4���Ta"yԷ̨�%=��:U��\�Ekz�^9�<�E�ց�"8�l:?��Y�??4PV�>M����Q$G�����W���`)�:v��pRH`ϣL'��{�>y0��`1��F�i��G'�:�0�Q�i���C��3�_���դ�B��G�d��><�On�D"������ �L�𤂣ʿ&�jm5��9��.�|�_��^���0�ѽgƪl����ݝ�����Yّ�b���U$Vӯ#�{�S��?+C>O��,R��hW��6����#b�,�ߗ��t�w��Sj���ΰ�ɽ�����XTLm?�9��u,G��Ɖ?L?��iV���IܢQ��Y�����LwX>��1,����:R�+��¿�+c�+�L����]ԚZ�Xf/��):�	���������g��K��ٳ)^DJ�5���B��%��>Q|(�'ۙ�)��k�<�qÜ߲p��<>Rۓ��� Q�c���&Coԓ"8�,fa �#�7�C��|�����!�9*�!�y����}�����c��	"y����=xZ4��"<>�Ԥ�Т`��@b��8�J��ר#~�&B��d@��<|���ib�.���=yz�dX=Z��*F��ca�6��f1w
�]��zT��q��S���y�f1��Ǔ6�n�(0^z���s�b�V��2�wW�Y�R
�\m�Md�K�QS�B
�|S�P9?H����Ӊ@�h�k�e�G
D��UF�}O&��H�S�LMN�G�����d�5F;���H�'4��!��m����.RX3��Mڶ~WG�ׇ�`���C�4xV��>�!"T��P�P��!�-\rJ��h6ۨ����A%�2M-���XZ_k�?�S4�,��S��-c,.d��nv,i�E��&Qky���>��Q$},3��MH�)ˎ�k�F�^����|�*^Y�����b&��O^�~���xt�Ay���L�/Ǳ��b�XF���Nc����i)�rƇ矾A�����x���.;n�KW���ϣL��W�����"2j�R�����4�K��{�?�� UzyY/ ^Y���\?}�6�'��f���	��=~��.vGQ��(}!�ʛ��Q���U�&Ɠ����HSr2Z��hC^���z7B��g:�6������ ����;���!ը�x.�ԍ/�*�����9h�%���CZ�H��#D[���B�i=yP��ϵ/Qv�P�j=6��<n��F\��c�8��\F�E��8 ��j��$}]d�Oh@q�0M��&2x�a�<Z��3��8��gvc:c}�B�28"������zn�����jw�7e������s�R�X�
eFׄք��R<�a^4���:b���G�v����Ќ���4��j��"���4e�Tk�T!]���,�R�V�sDyT턾*��:���Cé�=��j��ǛH�����!I��At=Q�@WX��0��j�h�Y8T�5�%��hWj�&~���6)��t��P�_B4����Y��M�Ē�	SHz�{��m*�.e��x�ݵ��ES�
mu�6��;��M|��,<�E�9�̎,�X�
���Um��v��wn��Q��m���G�����m�:�x��
Y���~J��r�=?m����_"�O�	�����U���F�V�A�(~$@9��2ʕ���1_V5Es�o����S\Z����+��8��M>`Zv�m��~�A:$��b��H��7�a�o��A:ٙ5(��"SZ�[�U�j����o�]��ܜ�+�Y�UӒ�X��:0�cڊ)Gv�?+�gz�(.��ڻ�ߞ,_���<�}�5Q�Ipi����3u�%��#�����#�*�^��so��X߆��E/�D��ǈ��ΡΠ��E7�D��@�B��[����jO����һ&�)��:���gѢ�nxi�gDF��ꉫ���5�J������A2��9�>PU�b����
:Ď>�|�V�\�x�q�@m�vQ)��-Ċ��R7�� ��n���:gG�(�����8��C�"�9�CD][��u�����������?��r���� ���7DH�J�-=¥h/��p�@ L@�Ր� �(��=̎��
 ¼y+��<8�X�B�K!��>�n<Fzl9���D�l�"]��S�����E'@/�E#��RtG?*�j��%xҋ?L���j��gh�X���B׀�u�3��4�`Do'J��d��I�Y��I�&xnm��Bډ���>f��Ͱ�xG;�;&pT��L�ן^�l6eS<tȽ���I��rXLF���e̯��EqL�v������e|�[_���T�>>��|}����?��W���~�Dw���9m!~��u��׿�7�B���'���4��3��o}_��+�]��Qu��U*�d����_y	�l�,`�>�ل *���F�Oū�?L�쥤U�okCTi�?�u5٩T��T�����C�L^jU�=y����<��I ����E��i�5
�2Z��40�'���.��@�V%p<�3�Ę�I���A3��jd	���F�s4�P��#���� ը2���Z�a4k�� ��q���y����zk�EO/���p��y��@M̦��� +��]�#3���w�^ی�8���Zu�%Z!MxO5M���n6q�.�"�
'i$Oh$��;�術	�>�r$�1xH�CZ������s>��w�ܽe���.5Ryя�.��a��>E�@<� �� ���\����(�%�M���1dy8��0��2>#4�R�Y�g��CD�x��c���0O�ʲh�r(ө9D
�m?��8Ft"��`[}���f��?��C�t�(����3�+X����NO�8:.cУ���Ċֵ��)ƔY�G4rw>�}�F��9x�k����=��
g;��u�7���ϞqWx=:�PO�(�ۜ`��j4��=ݧ���ǧ�|Ͼ���F�s����7�E�Ow"[��K�|��n(���j���XJy@X�E��\&�tR|����N,n�ӈ^Z̓��8��K���qk���p����ߺ���vx��j�l7��J]:,~�t�[ލ��D'�n�>�̣H�D}R�g0��1�Z�IS���%�	�)ң:Ү]�<Q�K�(o�L��[�$�d������L���[v���������������m��@�67ٟO����^���Ȁ9�n}��ګ�G��J*0n"^�Tk��;T��,��S�¡74J�1�b�4�����%�	��T�*iU��i��{DA��Xē`�p���R�,�<&� �aZ(���y^���Q)h�bT�H/��� �,C��[�F/�TC��_
v�G4x����³�����Q1�'"�:��|���@?xvϯ%wN1��wz~t�!�34
��͊��<IB2�P�w=�!�?5C�=�QP�ӑ��{����w}�|�2�gC`=�
RD_*x�Gߺ�_{��^�V��Q(�Y��z.�԰��l /__@!��l����3!�)�WGh:�z��s��IK#ީ"�s�����X����jЪa��g2�a�_�8N@���q�	*l�b*�Q�����c��Fi���]����N��8�r���G	dh���ֈ�Ns������9��u]��ȑ�nJ]�W�o��x��<V�iH�j��v�T\�$^�����x�^v�F�+�^�K��o���W�}�q6��ݣ���}�
~����|��|xR�L2����/��7� �r.������Џ�^��+�%hi�[8�F�5Hb@e�����>�hďvχ�'z�Q4	�����ݾN��� �M�!�O9	j1dMj΢��^�yTy�P���,�i�?D����f�tlE�	�o_;��(Z��K�O�+P�!�h�Y�)P2
�Y�rMѡ��)�9o�'�����N�<6�I���	�4�T�vҒ�RD��C:j�"��RN,����4�7�2�`�`s)���J�sA�ͅ�����חpi>�|pB�Ő|S����K`ZN��j��)a�MO�ZM�Z|U�Ң�Z��CP���o�i�k-n��i��M;2�t�0k�	���K��V����S�(D��q[�����%,�ø8.p��t#F>J�G;�!�@�t� T���M��m���[�7	�N�D��p:t\F�e�(iң�cR���&��L�k��Y�Պ	���3l�����8���_�Pg��\<,�h��f��1_���� ���i`Ҥ�e��`�7E/m'ͨ�����tW���
o�Λ�0���.��swq�����7��v�U�3��\qZ\���;*�ǣu����j
}W�t�����,gO�v��Y�#��߽��S�nh�`�&�]^�sQ�� � ���|�d>����)��%��7h�jg�۸0�̠������o�ۻ?�W��(_�u�e�s��S��h�*�.:�q��G������3n�'��|�0����4����"�����,s��f�	�ʀ�7@�5�%��a)gX:P�Q<���ni{z$��֯�o��9_w������&����?Q��wO�h�<w�i٥1���V���4P�I[{0C�q�����><���l#�)QQ��v��B~�~���ԗT]azE~� �&�Vs�/'c��F�F�������v��}2d�H� �ʺ?����D<  ��IDAT�!�����Mb7�S��z]�
K�`�n@�����M�x�2�$:*���m�٧/c�Jn&�e
�ū��q�
Vr�h��qL��_
�Gf�i�4��tp;�OI�ݪ%�Kx�#1���5��^���*W��h��-!Z�!�O����������"~�ۯ`ce����f!2��R�d��\s��o,������SX]_��G���Fc�kXnc@ �[YĄ�0@!m��|�(ܠ������s�|	����!C�V�II5ߪ���)�j�RHC�/ܧ�"m��&yc�/"@^��Ľ}�X���eTI�Z$�~���
J����Ǚ,������1��Bȑry��3�{U���{���,Ƒ���W�-��B��g�6�uq���sW��k_��k�yb5�?��/����4.�/Ѐ_�|��.��Qs��v����ū�ʍ�5������!>�i�b�?����<��8����v�A �_����Ek>S��o��0`޿�N���IR�vX濸U&��E@j�<�/� ��C���2%�:�k->�/S�U�4'�L��ݷ?���-顉f����g<�4� x �ݭ	�:��QAM?Ч�Kil��&"4r!-��Z��)孎�J��7��(�^[��?�������3[m^��d2�h�^���������o}W�\�>R�4f�v�2O ˴ET[�t���2�e��җ�2�Y���S���!�$��S�z<���F�I0YvR����k!X���x{����p�����0=������Y�EŻZ��;����gx��s�l$����n���Wp��*���HK��k+����B�<c6�'�E���KXZ��i���U�,�7�9P�)G�����m��Eg�&�=���,�c����a�Ņ��Țw"~����R��Mo��]�uŤ[���a�C���M�#�^D��{�x�"�y�FZU�2�Z�O�,�i���Э���~�C�F	 }��������;��Y�1y�=��i��$�x�>��,��{��s{�]��:Z�t-�L�) j�[��Qgqݰ���d������~�y<H���Ʒ����%��/�����4ׯ�c}m}�F.�1z��K,�%� ��,��D��7�7K��>����0��P>���S�O�|'�1;�m�pD�P��y�����(j{����р
9�cz?���I.�M�2�G<`j$@�����I��~���A�'j�6D�d�$?�D��j!I[�2+�|y�:�ڭ����"�����M����ΎO��b7���צD��ѝ�5"1�*��k�U����k"�m#ׯ"GᏍ|6P��$��a�W���L�tO���#�1��	��Iz�{�������<#8~�$���(,pU����iм*i���Z� ��Bm"N�
1�iTS�������T.ȯEiX�q�Sq������J�_F�v��-y1D����������X�{*�	������Gd��@��5e�1�vm"��(:�w��dH�\ J��l���MC�>'@%�?��/�l.�y�7"�c:��X��b�����T�'H�����q�zO=���*�TM����YXGq�^O�t�Q1ҠV��Nj�Q���n��J�O19}���6�.=>͙Bo_U�Z���9`��K ��!4}�q$��N�{'U�pIw��Sd~�F�ԃҳ����	L4tޓQd�ր�.����Pfᛝ!���R����ҙ��3� �'ETH���N��p�D[�E�ʮ�,��T��fm�j�I%4A�UAW�fȇg''6�@}�U�H٥���J�N�Q��SwXg�:n� ^��76z�6�,��Ύ��U�l���љ9�>_��:��5��4R�ߊ\ ��xTm�F&�����k�E��U�+3���>A�򰸋en1@,�B� -�Nb6�q�K�2�0R�j.��������;A����D�󸳋�������71C�J&�����ѡ�C`����w���f|�(=1�q�K@&O��吘7�ɣ��4K�C��Jτ��w�wg�pxgg�5:�c�NCay�J:�>&>�ut�Sn���5	s��v��]g3��Hc�Z3�t���!�'}�Ii���-ߑ @򿬊gt_�S�*-�-����#4���	����I�c��G� �S.�yV���!�:��0���9��!�!U?*-n5 �`�[e����t�<�~fn�$���z�@�6"�
|�:���h��՛�XҔ2����:�5u�6O�_�ߍ<G ��P���(���=,�1��f:4��t�[i|��Lݣ.�`������l�v�Zv�fw�.��IJm�e<<�o�p��HƮ�>���3��~�Q?8�r�n�����j����Gp��lg|�%��M�k�]�Y�!@{���S�o�DM_�����|zM��J�ZjN%`�������<�����q��
U�f��yac��hx %���!DI���[(~�>&:�I�Q�Fjv��w:71���HG:r�l�-���C:��������;��@^ �hZj&-­ZX�����_Tf�1j��m�%~�e#�Uw��-��u��w����^�Wf�N�d�����w�Cn_@M��7#8���,%m�2���v��P鑜C��1�{�ѥ�-U�i�&�DC����pu���kVS��� �
�q�Y�,!��1�u4:L�L�X�c~g���}�`Q�y��h�@�BԠgH[N�M�-��d:��%�>� (p�Xs>q!�z>f�Ok얋<VQ�P1�{h���$Ri��)p�*޾����1j����E���1�˝a�e�3�s��i�(=nmC�q��ϟ���X�W`Ч�I�G����4k�w*ݸ�@*���(����݇���6ʕ:ym(�tsT��P��,�����8k�nV�!x.����6P
�GO��Δ���}<D���Ƞ�A[�&�y��T8�βa�4ʚde�Hk����Ј#|���!=,w���;�!\�C�{�
��,��;�h��P}�l4w�ʼ�.�U��)e�4񩔇i�K��M���=�<�9Ż��p�����g��uk%$i���;���Q�z����):]>|x��>}��I�f����X&���2x��>���=���֬h��?;�e��[��`��1:Ud�=��y*�2���O�!��F�<9���9���s�7PMd��,J�S�ޓ��.�"� ^�gH�i�cK'�!'��,i$�,��bM�5�J�m �G�����+h��E����a~w��~�Ǫ%0K+P,/~�����D�D.�G.� h��i�����9��=��i(�4���{��]�d~Ɲ�Q�]����|�f� �����}�ޯ�C�Iqǈ�Jp��Y�0>�w�w7�q�B���qW"�!M L�`�]}�T����d��v ���k4��qV�ˈqpW��҂���5�ߚNh�5�n��8�p4�Z�B�	��KPSE�����<*���.yL�=��ffhD�[����}F�G'I�&DA��	��S:B���6�ȄF6A���<hɎ*u�P�9G�t,�A�3��X\��ѡj4���0jt�@�����2o�\d�ˢ�<�Y�=1�P`�C������Ae���
�]3Y�I�?ECݓ�j�|��� �i�y��#��.s��̶�k4�s���=���k�fdby�"���Kf��u�ٷU�|����l�2{wiM������3�c��$u�.�Z%��el��=ꇝ�N���:�6�(6V6�=�s{���㸨�X��X�N+�T�YV���-�-�}ai���C�aY���3.1�.5�K�ʀ@���`1��H-¯]����r3;�#�(�tW�`�T�v�?�w�����u�7��{�oۑqP����cRn����t�|~6;�c7�]�o:�Q塒������F7qSr�4:Ql#ϭ��<.�+O,{g@�z��}�wy����{��r�.:����w�S3 O��������c߳��0A�!�b\��>Ѱ� �V�N��֝!���JV!�AĬ!o�c�?�w詩��O�f'神�R��� �SU�c�>����T�|d^�F� �N��у�ЈQ�Ѩ;u	>轷��!��fpM#g:~�d���ҵ��&]�7�� Ul������q��WQ�L'fb�u�pƏ<Sy�R�'88��hKm8�\*�@,�&?�����XY�&���a;�T�Q��{�WC�]F��Ǘ�_G~f	���� ���^G8Aψeԏ�#%i���y�?n#��>�w�� �.��S�C,
B+G��_}	��(�y
?M�K{d���,%J��{�5A���tBP�# ����;T��W/��M�IE��+��v��я�2�<�^6������謏�ļtO��T��)��s� A*�i���98��#R<��l��߃�q��u4W�"Oj"�B'���y�i z�;�"�|�<sB^9J�`�xh$m�BjXb&��	�֟�W���&((!��Ȳlb�ʿ��A�Bxw٘�X��)�R�X�t��P����䔿�o��.�9���a*��0@��y���&���y�O������h����~,��썗�/}��"���<$Ljm�qhD��eH<h��љElK5��,r�(Z���4�!k?
��퐪Zʬ%Y,���<��J#.�)�O����Z��1�������p�	x�r4*������tVri��[�'}?NV.b�[����=�W)G��~�1�Θ���j?-h�T7�K���i��py��C2�"O򽩼�2_�%Y����ja��9B��S�9���F�X��=l�p�n��Ѡ���Θz�V� ���O��m< ��R����s+�V#9�[���,�w��&�A�щ/���U�f.�`����K����}:R�dl�����1�n2f��Q��9�!�1��9䳀� X��N���Q��r&=�۴���:�ّ\�F��FRh�H�gz������;�D�Y��=K����i�u�Gy_θ�14�J�u�i��i�$M��k�m�|O��.�]��w� � ���L� �;X��Q�v-�/N��bs�U��m��Zҋ����.�_<8�;�(�D��¤�`<��J��6_�Sܥi ��Z���5��"�#+]x�ZS��QD([!r�j	���48By�Q��-e��>�H6�R��)Ϥ�y�ժ�S�"����B�-?\��_�ū�9d��6$��w� �����mv�{��n
�O�8?+i�?���wk�t��w��������@Ӭ�Ǧ��%K����Y0}����c|Zl��C$�5jw0��:���&���s����җ�\z��h�N�1A?�h�:=7Fy&b�����RrQS��dh�.uNմV�X-���0&�.I ��E�b�<02���AMqЮ�E�w���E�=�S�[M��L�O�5��[����*�)2V�C��oz�ib~�g3�2%"��Md㩪WIpK�)%�M�+]J��M��KNR9��|�0���D}TԷ,I��%=��4���0��A��k�/\�װ�!��h�|e�*�`(�v"�����:|ҥ��$"�+/�F7@��ma��� ��O1iU�O��+�>�M�����ǰE�V�h}j�`z��li9��]|�� ��!�l7N%[#�Un��f�nM��{R��FDC�D��6�g.khdbx*#�}!�"�i7^#&���5�_�G��&��O`���(��Ry�yt���e��\5vkLw^� ��?�5/�9ܶN� ���@�X���8�.���z&�)�,o�F��9�9���4����-d0�DC�	"@��o�d��-���5k�8C`n#��'&H����T�>eN0�~܏ y;�����a��ѧ�DBL;n��F�x��`r|���Q���Ư~�l6����
�K$2��ٵ���!�ä�ktU�d`��uB�C�Ox�N��!A�Ǘ�����R��Xy�<i��LTK���L�j�� Q�$��ir�	��C�?��LKǗ@��e-vH�%��rD�^��i%3,,�YX����n�w~ANifri��k�k|r� �$E#�xP'/@M�	�ff�DR>Ϋ:���и�ܮ�k�gm����ǰ��&{�L�,$��L��h����Hh��C�	�j�9�|�%����򙁺`v���h��e�6)��a������L聙5xV^"k��1*`8������i��>N���O#�j�����m�t���Ƙ*�R;5��@�8E`D~7���Z'O��@�K�Xۈ�%�j�5��묻�ݦ38���ae�k;�J�� �]g���\D�k��5A�t�� ���Ӽпɾ���xC����>5�t2}���/��7I"�ūjo�:R��s���[t�N��z�w�o�?[��h�=�������-�~p��"i��dh`���	ѩ+�Bp�N����`�n�����h_�6Fk/36HKs�H%?�����;�Ai��4��)�87�v7O�תT8Ͼ��X^zwR�)�u���a���: 3V�2a�>�]3��(pl�GtV锻���f$���[5=��硾��QV%#a��F2���o���y��*}znN�F��O��wD#S�EE�-,c��S�̬�Pf0��L{���Tb,X)eInyZRZ��B⹫�X@|�vn%c�5�υ�8��B�KA0ŭ��`᫪^�G��y��L��l��R��#�/N%�����4�G��R�u�IE(�1��ОP�В1N����.����)!"�v7Yf ϋʀ �$��_�g,��b�ޤ,�'7W�%)C�J4EC����F�nO��4<�y
Y��k� ���hV�	Ѐi�h�
�ϼ��Z��+G3+Ӏ�I�Ge��W'PhL��hskEAz���<�I|�4����	���A�W~4\]#�tQ�� �i&�ճfZ��c8��~8 6�S�U��rV��y�ʾ��]��֯B����<���=�]��*{��i��)[џ�!/��F��O�)�l�>4l\ob��0P>N�	h^����U�~��JG3�G	0�Cz�Z�uL�L�T�=5)?'Ux�U�J*h}F��ƹ4D �c����eh�P5��y��!0v>�&#�9s(��C��	Ԣфz��A~�vVM�}�9HXB�i���{D��.|w-n��ğ}��+�'�XY�E�P@�;��oW͉�(�K�$嬓+7%E��l��B��#��<�@yQ�LuÄ�E����f=:30	�)k�E9D4��S�urv�$��4	�ԏe��*to�����[�2��:��d2�Yr�feq������;��!:��x�ݤ�� ,�@��1J�&o"ɲ�<ɓ�{��K�&]��w��wʬGS�P��&b]������:C�|�=���� ��3���,�.�4�ՀQ�yD�2�1L�0`Ւ�ttv�!�4Z{c��a㻑��ٴ�EX6~�y�$�)t�i��s�e��W,_�!�-�5`ِ�>�t��������t���?�O�u;��W�'�f��V0B�r�T:`v���]]0�c�������n1"����(����)<��uW�t�0C�^�[߱<0���<jF�@�a�[ԅ��Qn�i��I���1��y�6-� ն�(���,���~o�e�p8���4Q��x��@T��4�s�õoa��J�"�k��W�Xؚ�M��ԛn7҉�j1P>��i����ʾ�)�K�����Ș`e����������څ9k���� ��Q��"��py@��>�,8/���{����s�����~9��� j�3V翈���7O���o���*
I?�Ԑ��AF�U���� �/��bX�� �j

�N��	�2->��`2�Y��
U[�6�j)��U�l�A���X��:��T�s��}S��3�y(ba�=�U�Z�R8*"@P�M�㣱tZ}}��ӣI/�?��R�U�3�������Es�6wsYN���o��U�k�=n��P@��-0�Eb����{�ie�P^c�ӣ~�(i#��~w�D[�¯>

�H՘�\^��e�a>|ҥTZC�O����q2��,&T������k ��K�#�xOSM3.�T�GT�d����o��ĸ	�q��P�j�z-�3�hT��4'f҄��W]:)*s�P��vL(�,[��h�r�7$r�=##��)[��	0��Ji�-��r�;��~(A;��`m�ت���f���� �F�����v�2@�|���l�:C�.b��9y����s�4=����e�I#i��Fk]�������+�@��O���)�7��P)�g��:��8�����ow5M���Q9RAj� ����5'N��l5tD^,� F-�d:a	
˹M қ��0��¼8���=)��"e':�hlmMM>��*�ut�Ui�"aHC&��`]�o���?�a��*�;������4��gii�a��T;�����G���'%_S�)n|G)�7�'�@��Ep�Ѫ�(�kK4R1����(˲��"1���,����o6Ѓ1�����0:��m��վ�zVH��'R�+r����F�y��e*l�Q8j����>9�t��g�ZLs�S�r�\��1�=�iF�ӳ��t�&D�#��z�+E�GzY��|ɡ�������ON�J�pL6��)ի��I#�KK�B5Q"7�_���#,�\�t�y	�����sZ�Tr�w�l�M�D�YD&�v%;��5~�|�"{��D	2��{��mB�~��V�����1:9}��dX^���[�t�&*[��9��1�3;�d�������ń�M����g�壹�DW`�c0��:>wz����ȨMpݵ�@�xɕ4E�5F�2��i}�6����S� �ʄ���5��͖�bZ�Gӣ��Q:*>�Y�^2��_FC!ɌxBd	I�MAT��.x��Q_�8O����PK�Pm������/ꝃ�Q���S�)�����{vt�����M4�#KjB�%��e�7���߽v��gQ$����1��3,��C�� ��zz�Ѐ���ƚ��GC�h؄��r�z���)�.����@JD���j�u`��LZ�8�s����J�I$:�����Q-��dޢ�Ũ���$N�pt�x��!C�
�A�B��2��C�o��D���q�,�W��ƛ���NZ�K1_u�)���<Z8�j�V~e$	���⠌�:�RqZ͔��HFL�+����Q��j��d��;G�U�cs0ɀd	��4Q3�sGs�"A���������g9�`�S�Ј��A4y&Az�oeA�1num�)�]�Q�Y��cEa}ۘi�h|_��q(>���J!q�6[9� �p�D�*S��R޺�㟂1�VFuї<��+^�����	`v�P��if��l���\t4#�r����6�fۚY��c��aP�1Ӻ�����'=EM�H���_���S�� ��&m��r��z��E`�!˱�<��'Y�ZN����į���z��$��0`���<|K���t���#�T�C��Go��<��,[*yO����>�H��R*]r������ъ�#���뤁N%���Fl|����1u�� F�k��n�F^�����͹�F&?�����8��#�:g'𝕨�	 �A��/�y�x�[4�E��H"�xB��s>�m�婦;�����xCt�7�\/O�ra�i������ZE(���+��V�tW��%��j�������(I��`s�V��:���q�Y�j��	�j+ERB����~�c-נLPZm����t��N�$�����V�gZΩC�j��4�Gra��"�)�mf��	�ɗ[��I{ގ5��@L��jC�>������j�U$c�K%d�T��"���q���Z�U5�2.�!�<��:a�\��q�3��]�a��=�kR7��oI�����N�xaFy-�e��f�1j9�&>�;��CTB�4�j:��&��c�'9>ʻ@�'(��A��B��Ͳ�0`���VH3�!�C�����Lw�2��e�M�fy���}TԤ����"`R7@��C�<wB�툸���O�jhD%��0!�::��&�e�W�/2#b<�C���-����ե ~�r�ݘA�@M��G�S:gT�|��bX�Ho
����d�:�`^���L��6����
Ǖ�_&��{��Sb]�����My'�$Ҽ�!gAq�o���V%�|�wH*S/��Ǔ��N���w"���~OS�V��P	֚pju��D�*F尀�Dge!�"�NE� RLjr��`UK�JT2'ap%E��wL�z2�@�����D�D�7f�`�[��C�a��a�Vq��o
Mτ�y�>l�o�k�
�H�~�O��\
�	exw��O��B����ӵFY�{~O#-�>M���2Rª����*�1�qT��z!��k��!��qPy�� �Z��vk�Di
���.�ղ7����+�!��*cM�)/K��WT`�>x̣�+���Y�
3U��6+0y��T��O cs��hdh�a+�9E���s�a�j��Nu�o(�N�`FR��5I��+�}4�6S�2#����t�r�Hw�@��� HQ�IM3 0�f�'��ۺ�c<�q\��FM�&MJ2�0Dy`>�X#�
PqNԼ)�N���7�Mh�9f��h�$���ߵu�������yd�=�A�Ï	�����^�Gi��]��-E�c�E �@j]���֔5�1-~b�l�l��95;)-h�B�2��.�f9�lϢ�@��+���L�J���H��M�x��uj�\	�[͍��/�d��ԌɰjZsT�,�%O����h8�M��p��W�+��'��Z'���cĤ�A#����-�T��te�a���F���(���<�.�R��\Y�]+��uOv.�H��P�0�|��Cn��G5~��#M
k5�����ݳx��J�	��ԙvZz�:4`�|˘Ӏ���"�Ъ%L�Ӓ0�eM�9����<Z�Y;u2�LZ*�g,� B�2��R�=0],_ɽǜ7ɲ�,Z��L����j<5�L�����WS^:e5Ϫ�R�-n�Q�P�c��G+gm.-t0��3��s��gn9���a�©�t��yi�y�}�ٮv��:���T%A5��Ko�����	�5��bvlZ:��Y�@��,�,���#2C�=���k�W�)���,�9�4P���D���SxU9��UW�T�8�I�4]ȝ�f,�*���&jRd����u�Q�X�m�W�*ٓ-P��\����d W�\ʐȱ"�*��'ŋ|�*4�m���q/L2��dJ�Ol��x߈鞟��%l��k��=�Q%i:����������&��?�ƽ*�
QvMm�F.Q�a�j���I���>�[ۤdA)SF<Rm�IC��捩@�<�0��M��H�#u�z��S�O�P�y44�w�dZkMl
��$R�-GC��H�)X~S��z]� ����Ѡ1f���2����w�Z?)},~WGfߔ��|ә(l��y�$�t��0��8D8��pf�]&�\b�~��"�S����&�t$!d��'�6��2V'P�����J���H/5��Sy�i��� ���T|ݶ�)�H�<�48�uX}�c�/�u�a�T�L�uY~Z��d�2!,� ΐ`{�݀����_+/�m����|�K�}�Qg��"�Z�c�֔b��7�}*� �_t8�-�W�X����=�Γ��f��_>�:	�qS+�G4���󈚸�$�=M�  ��5Co!K�"�t�5gћ��/�B6�8��H�(�*��LL4`���7�g�����eИ�����!�z��b��S�d5DI3�u�c�O*�H�yy��,�0��4�������f�C�?���f�:O�tQ��Ey����J��>��HC��``X9�S)Q'���� ��F��s3f/0F�����*ʣ���ɬ�;��\���H	�I�'t�Fh�Ԕ�)�.2c�/c��z`R�2�3YB{X���K���J�(p��rl���܄2=&��UaɔӴ1~#}˴?�Y)� ��6]�MɎ�I��ӹt��ƽ^!��|A�TӬMr����{n�r�$ת�s�h�x�;�S�I�Ms_�H�ߨI�7ɇ�L��D�����<�+���:N��{�!NQiv��&C�;�R������t
��F�����>��4��ՖQ6�T��#h �7G�6u�/p�����7ՇM}M�k�7���@�H,�� +���UԼf�f����s��s����ª������6#���������M�+�#�M�d�"a8�?O����X�ך��� ��!eK=7P-���.~2:�JOh缪��,)/G<*N�`�C��"3�:��~$��ߋ�Ȓ��pWl�#�m�y�2�N�ʱ��(�hg�0�%1𨂃9"M4��N~�G�w�{�C|w)�߻����t��h0�F�Y���T�-v}�x�b1j�4<�'�)����ܦ�
��&�Q,l2���,������6����aY�	�Kޢ���� ���C!OSq-5q�i �-bw���z7���D��v��:�B�6w��`gSs�ae.�D"����)4�i*� �4�4n�T��C�[��T(Z�#�L��X�K����)�(�&�?H�LK2��	�z�����	Xɐ�:b�5��*	�ΗR�M�L$2r>�=&�~����#�H#;��.��7x�b�&��)r��K���F�H���\ek���ߍD�*E�r��biP�d,�g6Q �:���Qw�`ЃLZ�2�~�ߢW��8.P�^^��3>��[�}�)\��������N��?D�Wv�}��>E��A2�$()�`Eћ@C��*�L�|���m�w� N�dyR�$Ĩ���,�ZgW�����}�g�i�."�P�P�h�i�E�S���V��jBxA�<Rqz�uA��I�N`����4���i��:�3��'j?�C��w�X�qe	�r��˞���,z��D�И�Ȃ����3x�%��|��a�tmLY\Ac>N'�Ụ7���$�rV���r�Q�q9�G���n�(�(����ѧ,h���0PM/`�~�j�4{���}8I*`>��޽d�`/��X���9�&�$}V����g�G27KZE	 H�z��G���;�0�#�a8�A'Ŧ7���3�$,K�6��Kdy��[6�_�40�{�]�(�&]���e�N�k�n� ��*��*n�#���`�J�Int��^m#ic��j��VC��E�3�K����<{�L��z�'/���џj%5hb(�N�`\V�|�,��w��@�2���:��s�r%�X�(�ld}S:����ת%P�v�[���F�O}��.�Q��{E\�Ԑ.n#Dlie7��b��2�9�b��z��hc� �^��`�trC�4*��d�`�Ep)�A�A_`�_���<���
���*��>u�� {�ڏ�Z*j���
�y��qzΕѣ��:�L4�]���D��L�j���v�.e�>-�sxnxe�D�>D���E�wn�>��}N'�N�K�M��M��E��Lһ�߂�2d�d^��4U��Z<B�!�iv�Ta��'�F�K-@`6�q!j���>�2�@Mt�x���2݃�4�bqiI�a8����Kx�@��Wg��;>���a��x�9Fsv�ܚ�K��$ �Q�/��t''J�F��b�w� jc:;C>2��y�p�o��t;��6�N�FF]L7�~����h�-�".%��R�����/B�츃��@TI �/P��Ob4^O<8�FT��ZϢ�߼���;�>�eL2��Y�F/7�������q�&|x@u��CPT��`&J�~'���S(�f$�y��)q��=$��HO��D<4Y��8��L�%D�E�ɓ�5p�ӀV�G$���E����
���Z6��оJ^ C��j˔?4fP�"=�:ν~r�2�3�Pq��O	,��W��ʂ�:r���P���Ui�^�.@$Q���h��!��t������L�M�(����B��r#I�q����Ы�q���l ��o��_:�'���/Mᾎ��7��B����T@�8+����;8ܹ��{wiDf�Y|܉bk�B1��Q�J��]�.Z�+X�G�� 3�&�B��!�O�Ґ��+�5�̣��E�z�Z��vl��K$U[�>1��u�!�L���5 4ڞJ�<�	����r�-�=˪�*)���w*1*EO\sr�ji�� ���F'L�P�d�X��3��.���#��$�uLJgp�4*� B�. ���:x���@<�G�G�8��0����7�
Q?�G�p�e�4��e��	�\?��̐�[-/*���BI��c���� ���FP0��^ď\��7��ͼ��>��
��$Vn\�ƥ��BZ�:�>�}���n�sv�����!z�,>�F�~�2��%��;�
�4*H쾅����f���ǽ���s�N�]O�'�\�~�2)�J'�j�%�7n`D��6]�6�ZW�?}��2ff�լH2JAk�k^��q���D�sՌ�L��-�fܮ�� �&�)�򓅜ʲ���L�qgxɓ69%��<�定8�BH��ט&�}^��n��rpܾ��֩|N��b�z�d���Q���N ������L:�x�:�{�[�J�f�V�\�йi�N��4�{�}���O�N�ǟ���㌺v2�� �W�t�1��|����X�q�Ƴ�11�Jc͉�m#z|��K���5�'-���6��Z׿���ŋ%%��\�4%H�)���@ODM��Ł(�R���"E�@yw��J����.�o�x>��Žz� ����8u�3�=�ta��a���`�rxi͜T�]����3�~'���]4����rx�ŗ��fMf�Hϒ,,�D��Y�tQiWq����|�#�CI���wp2�\z�ȭ�+-�#�=��{��(��/�񻗲�Ս�	����,љe�5 ���Ol�d�A�12>D��<ߌ�<��	�x�@�B֌%0@J���a���|VeU���.E�*f�y����3��?{uϬ&q��oUĩ�4"q[����]5�-z�]�͓�����7�@�>��A?�Ϡ�[A`���SCj����;���WfS�f��Ϳ��{�����������ve�\�����D"�44���M�Y�F�y	�Un�%�
XJ��{�F��t���Dqؙh����\	6�Zm�6�;�j��={E�k1<���Z_�����k���^���_�@�q���w�a��V^j��ȧH؇x�+�Z��C���F�i����5xz��^�����HƆ8޻�d<�Df�8�?�/�{X��L�"(��5��_�9���U	��v'ɋpRs�|#o(p����~�r�.&��a|���8.U��v�)�����kX_��O>z�Zw{)<Hm����8B��g�m5�)�6�S��1�*��i���h�4	��Y`&�Q,h� ��Uۘ�U1����0i�>A��7�pk�FA�˧1" P�(+�8����S�^�:w�<�����8.j A$�wZtȃ�-g㋳����=��>�3��W���ek������~���tL���>��gi�"9�K��W��6��;�=)�5����n��G/��pv�NW��/�q_Zϲ�K�:T�1��9D���K/�|땨������<�Z	^>y_,�7+^����s����Q�. F ���.~�jsL�����_�G�� F��f��F�[����"n}�N:q�t����*��O�H��Ź.}��BSY�Ù1)�]-�"#��òVS���5j�RpMO"wQ�gN���ʧ`�j}�k�d�d��ð&���6���o��k��]��s��W`BG�������];!ߪNN7˶�ǰ�J�p�C�}��\L����X�TPm����ai~򋾦����&Mn��8���w?x���$�;���I���F~�P�������na�W�/\_C���:޿}��5�u�o4�s/���k8����S������Q_�Ng�@N5��U�W�2~�HS޸db��&�S���DIo*�\��37s�tO��W�����i\o I�:gx����A���r,�+��GMd����g���%,o,ѱ��;9�?{G��q�TG����u�c���ן�V?�G��9����&ґ\��?����F�;�$�Gq��c\~:	����AUgZ[�Y�a����ۿ!��(vc�����n�
<W��1��!?�V��@�����@������9|�6�4�(&�x�$�jyE#��9��[�۹KF77o�sm�������q8E�Kھ���������FD�k���5�靻o�WƉ���W�����xjx&;��kY�Py�R!?�T��P�q�2^-V)�	���!KҀt�-*x1��R[N}z��X�L���5D���o>�ǟ|�<��,.�#��<B*�7��e\(�jr��pau_y�i���⣽"�Ԅ��δ��C��#�%�|h'Pr�]�*d���4d�$�|n�rw�W��F|Y������D%�J����K�h��_��ՙݭ���1u���'թ4�>��r�ڔ�<��
+e�8lX<�5o�|�3��e^�4�Tڈ�h�g����L��]��%���x1�ŷn�Y�|2�fyh���4\"��S�����A'Z�-�@4��G��7B�ԛ �a�;$m<�����/���\���
�N�j����,,���^\���%U��ePn��+ѳD�'��ؘQ�����1�vi�<Ѥ��ۧѭu�H҆��C��i�6��5�&�q.	o� ��;�$�������T,��W�P;x���Xo��/������	��`\���]�7T�_j�q!Of�py�u\���W_����ڳXՌ���G�����6V\ݸ��^xK�����ťIo�Vp6���jĬ�$�?���g1��;����W���G��/ᷙ��5(0䥢f�{�mb��z��۟�;�#33����6�6�vz����5jw1���������W���N��NP-\p��˔ӧ�>G6�ó4�n�#aqf�{%R��%xԷJ,�Y<,�W���y����
?D��%�Q<��U�E�}�A=�Dvjj�A��wk���ϵ�n����w<�τ�R#c5HA�m'XШ���|�:��6��Q���4�F�&<����#!��I�������g�Cpܧ��[�?�L;���	�5Icl����8���\\_C"1���#�d�դ��N)Ķ����&8�H��8���U��q���Kt"i:"�g�iA~���,���^�+/=�h6�b�%򠏴|��Uܼ�&��|��4��]$6���*���>�,��Qٙ�69|���O���-����R��6���ṅן��O I�@��#<�g܌�������mv���5�m�L�(�;��Q����k��2�.\����\/�ը��<CP�&V�Z]{�:��.��0��̲���
��a��>��2r��7���ʳWQ�]�Lh2e����V�
\}���>��QuU�R�k�p,�L!��J��M&�]@H��L��N�a�;��s0�⪕��j0=��FB�6>	�ޓ��>7���Q��p�{�>ӹ�r��:ک�𡅳���m�5���ͱ�i�;]^��{����:��Y�AP�'�h#�0��+���a��x�|H�2��u�H�!�E�ĕ��q��M$�� ��s豠��՟!�8������SU}T��89>���)�*UTk-
����~�.��,0-T��D�OR��ȝ/X���eT�yc���Q�j�&�'�X�T�3����H2*���ڧ;��ٝtQ�ow�YT�Z��G	������pZ�ԝ]��.�Ͼ�����<5�X�A�ϣj�,n!!��n�?�ݎ�|N������h���Yrdl1�:?h��F!���Z�1��Ma���:T�����a�d�@��S}��<�W�c^5d�ϴY�.�C3��?AWI�l�����95�8;8��[w���j���6uR+k��t�2f�ih�Q4e��	4))��Q�X5P4r=�'��i��4��c8�t3o�iQ�T��� ]���jr���_T�C�,z�>*--	䉇mY!O����!`���I���q&�a!E��=�vL����Vj`4��-���qI��14zc�V�����I�C�v��"v��q @�Z�P�&j�������MC>���<����;P��r��_���� ������@��Yq��L�<Ȓgqb5,��|�y,�����s!c�L��5�Q<B��S@��!H�Ndr�?�{ՙVS1��X̮m ���&�TS��I�����+ͼ'~�l� �h&%��`Y�	�����X�o�v��?�pq���]��8ȋ6:���1nuR��H�l��gGʻ�|�d��o;u �U�F����E�V�����шQ��ʌ�L�o�����[����'���c��SAʭ�@sG��H"��4:m�XF�쮏��A�&���&u<����p��Ud��G~��4����@J#T�̜���a@C?��~�j�.ڌSMj�h� ���Y>����ҍf,�dE�2���n0�J����&0�o�3������k�N��[+�w�=:?�����Nܣ�ө{���O�=ҹ6���R�=��4� ��G'2@Nל��R	��4��tL�h�]uh�2�\ܘ�|!I�< �����t���!�"�g��.�/��1n�%gb� )�C��_f�I�KWo��(d�}�o��C��$(o�;�gJe�6RS88�$��9�l���d��`���mk�3��l�'���?����D)s�01�+�S'��o�W[Ӛ(����9�$/$�/E���N��F�У��풷2���{hdV�	��;t��M#r��s�rgQ����NM�X���;~zu̴KX��ax5�m���n���O�m���8)#�G����~ǃ{���G%%p�}�ʊ�e&�"C�bS�R�L�+�Rp��[�F������9����bX7��辅U������K��[U�s�����Fn)nn�~���=���$
�v�T��g����h�T)n�GM�dD�0 ��K��j��w�9uB�:�)����&��;ۤA��ސj�~�$5�|�]�mx3�z6����<��;8�vP���s�F�y�����RA]��{[���~���[ح�J�ԫF�%�X_�@$���N��i�H�|�c~�=�� �<'gp5�	\͇zp�4Z��C�M�b>E9Uרht�j�-Ƞ�_My�(�h0�	�TOCѦJ�so�^7�O�}2����q>(�H'���|�����,Ǿ��� ?�,���b��� N���7�������y�6��$@�p��_��ƃ�=,-α<r��<¿��/pzX&/�\\ø0�a(j3�k��g��<:���y,�b��Э����	����n)U��
���e7�� �!A��sw���N���'��y3��]F����ӪcԨ�x������G����Z�!��sT�9��3�oo~x��%�VAP��U٪\xbs�� %��z���Є�1\�r(~V�|[-��cȫ:�sɯܠ9|4}�X��J�������uϦ��>2�����▎bk�U��Q! ��:1������www�c��<�IG���cO�9�hc^���0���R&�W.� :��^>���C�|�	��Yf�����4.L�j4�[�����x�e��c�g9MJe��I��`R�B��%��츃;['8��p����"f�ϹX��,�3:�����[5t��!e_Γ9~�ҋ�pS�&r�;�k�9�W&���+w�W�k�S��7-�i�n��a\����I/Z7~E�w�]�I�����Y��h�a>�A��p�(���XW�wno�/?��;�u�/[=̧��3d�>�`o}��{��S�S�+yzL��yGxa>������ʵ2���ԣ�|�,�[M�Q�.�%����6i"E;E����|�gꛘϒ	�n-;u�2!9��'�����J.�+�'ɸZ5XJt�d��1�������(
N㚆��Q�szj4�8~��
���td-�h�3��6��x��J_��D�f����5����b�"�T�^�����l6��h�h�e��D�~5qаkr�(c�o�;�"�c�R��{E�"��8�g'��{x���G(�k���h�Vp�Y���UTӳj$A��Gk�Cm�����?~�6�Dћ�HO8�fZf��(�*9G�F:w�	����T_��
�h�]��&��T�H��(�3��)~k*S<�wrԉ]S0���8�f���Q5VznM��7܉����nե���}K��M�ogJ���>�j��2����X��ꛆ\͑���Xxp5����'x�ћX_�#I��#0�5��32�ѣ�<UG�A����!�s��ǝ[��-7P�L#9����i �=��A�������}�ŝ}.Ҩ���ypX��� ,�Σ�����y84�4�R1�W�|B�h�쨓���S�@-`�LR�������!� ��t$��%j*�,@��c��u�gMCI�A>��:��v�IGh/q�� A�f�����RG�Q,�8�6	�3$-h\Ֆ*���qR-���^��G{���';��Oc/y;�5<lxp���[1��s��_��C|\u�[���(x��N�8r�_`�WC�w��-g��p�ӷѫ����P&��{]�]�&k�e��N�e�j�r��=x�����c��|7B����GpL����6��!��N�d�7��g�w�l�r���P�Q=)��3�1��߾�w�-����y�a ͇$@b��ȝp�`G#�4L��rM�b�E�!P h�4
*�Ƅ��4NX�C�q&'E�=G��4�BC�0�M�:�I!����e�\t||���'ݝ�m�%�e��yƗ�uN�R|��G:2MN:i����J'��X�4�i��=��x�s$���A>�^!��I���z��!S?1p|�Ug��b	M^�[m4OO1,��	:��eҪO~��}�ww鈄�I�^Q��k�pwo���#DgVQjD���6~��`'�<�j=��?�O��o����g�g8�S�G�T8�,զ���&gNJR������D�G��cp�3#��ӝ���龄Ս��u��|f��+��~Sմ��=�c���i<���+����{��l[��a��s����z�U��]���n � 3�f8C����A��qH}QH���#�I�(C�H9ΐ3�c��i��������=��~+���V�� @�y�>{�4+W�\.s�Ν���W7:��r���z���x��oǛo�o�ދ߾;��d�X�/|6vZ�7��Ql�W�[g�_��oėc��M�]';���t��n\�3 ٻ�o��v�쥫�s=�<ފw�1w�i;}���%|��<���=)��|�i�ï�;�e�(dH�"���i��צ�&mJ���z+>y��Nݠ�J����Kp��IBy��Y�J+�F���,����ɚ���ɩ����>�i'���唻�ʐp5*��q���=x/ܿ�^�>5�铭ئ�w�z�Q؇v���>#�1�}��SF��/��a|��Q-��V7��Q��O�4p�Fq��Ӹ�?���N|��~��S�'�^���Wc�v:������#���o�η�[[Gqp�ň�����s�c��[b�ڞ�;�Ԁ�qi� ]���)�M�Y,T�(��a	�SF��'Kx_��̌��.���$1
�;s���E��)�!,Ҫ�t��w��(�e6B�>�-�w�;�	�Σ�q��E&��]S2��� zOލ[��r<D�>w�f���<o?�Ǉ����(�=َ7�|<��Xz��2��G��ͯߊ�r}��-��oJ�X��,8k�{���v��Q8����q|�G��͈+�Ĵ{&q����l{�N�N�׀wt�zDg��Ds��a�߾��*Ֆu�:��O'�v�\L0P.��1(p�-����,1�{F+���|]c�,�m�w����nu{i(�;۹����t������~��������<SW��`l���f(Ή�\ϕN4��=�qFv�ވ-���qp�^|=���c��A�`�оo�݋o<�X^}9�7^��n�C8'��#j�-�z�`+���E���֯���Xټw��[o�?���8���������1<܏��v<~�omů�w?g��^��7f~*���޻�4C�'K�⫏G��~���1\�O�;��}GS㗿y+�]��U�8>FT��&��`a\�h�}\��t����upB}t�3R�p.�)x�O��'�Z1^����'�0�n���d��'s_����E��|}#k	�9���e��Y�ɣWg ��Ͻ���_��8�h�Z�T��pa�fz8���{�L���g����=���n��y��׼�p+�<xw��7qn��ჸ�`�Ç���7���N<�z������p;����]�w�\�wV��t	'�y�h?����۸�~<��=ƭ�+qp����b U�,�E��N��n?�� ��?3x4ߒu�4d)gʝ�È�	)�\�������xO�+��O���JL����1��!��*_�s,���6�.N�\;p�➳Tu!����wS�N��l`�Vr�����ߍ;�;87{�����M���s��19�bb%���i��W�k���;�bޟ\�T�<b�����;5��3���	5���;[�%��~�Q����� �x��w��z����>i������q�~�A�Y�#pgϠ�DөʳtA7`�_Xo�Du�	��l[O'�<)���,O��� $��,m�ş'�/�0-��������|������F�a:�������jG0�'L��fo_��)-��՝[qax/�MP���#�F�\�i���F4}��^8��n�3��@ �{;#��(�`F꨻���L�Ğ�oEG��452?�˞�`4�0��~t=������q��'�0ԅ�����NQ�9�P�����4J2�\ΜeWs�F�jM�W���9�N��S��P�s��U�4�\'�ҁ�5�͐�dc��#7��"c���Y�d0��c����8�kC*�E妧��4L9�׮MS9�GQ�7�f��/5c�uVl+O��ٻ�K������8�{���،˅�ӣ�ػ�a�w���s8����;���ͥx�y&��n�V�i�<��l���FL᝕�^���1���OE^_��XD����~tN-eێ4W.���UP�q{���t+�;����a|�G���c�'��Bs���I#qzN�p-ͼ�������NN����֣h�y�L7����l<���{r�t�Wp&���c0�qnE-�W�}�Qc���ݥ�<�����T{-1��5F�(m_�?B�Nh��Rf�&�h�����²�\ _?	�a�@�����;�w��v�c|��~��h~�O?�ׯ������{ă��Ѥ�ڧN��(�ѓ'���"F?�㠵wG�����z4NUo:Ⱘ�'�a��j#���v�1��j��E�j��1{�AtF{��r��м��z̆�t���Gܳ�"О^R���?\|p�빴u���jL�`����}|�li�1mC�������G�q<���Be�*���>�*�.��*�ǡ�u�����mr+��kF-@՟sʦ��}�|/N�h2�l>�0N�ߏ�W��x<(����J���mx�=��t��hn?����X_^�Y�[&�/��u	�𻳶>jt�~��`����h`���a����z�R����>@O�|�l��O(M�725��[��>J��;u�|ʭmu�X�q�N�S�c$�4L]�t�ڪS�p.�HZg5���A�Q�J$�T��Sn���R�Kӝ�������1%�����s�?(�g�r1���h]�����8h�4"�@�Y�_�Out���7M�N������O�҅Sq�ӟ���;w�=�}�,�ve%��ޏ���X���6�r��	����X��ƅ�����/?e���;�4i��I���n�͗6�/�8ˤM}����p���e��8����q2�5ϴgAÓ�~�^��w2��;Q������RUX_����_z/��sA*J��n͏2É�E�2�C
B�4;<��x?Z�j�({��{�L�҉�vɛ���E���<�'XF�~����;�jW����H?�� `��L:��ߚhS�h�̳��0��xC�i�6�~�|��71
�(�>��H���2@�\�D]�H��{<�nP(-P��aRla	�{��m�N)��HG�5�E��sa_�w�L����CQ�*2s���+�lK^X���m'CAG<l�$Z�Fr��{#O7q�\�[�َe��J+��1٦�O]���+�_E�O0h8�{w#�GXwQ2������ڦ���x��]y'���R\S�F�7yt(p4
��'w� �	�qhQ�{G��>w-w��=�xt��`(E�����"N^����j����5^b�O��4��J�e��3�8��-���8o}��"G�8���=��i��uh���b}5F7���8|�:��4�@6��Y�{�Q��}P�0��>:�γO}�?7|����^v�}'�-��6�q�����Ʊ�<��p�p�\�ڂ(�.F#��e��8ak�m��PV"� �	s�2�g�0��pL5�\7Z8P���#��1�f��n��'��k�&u�Fv4���R/毽���@�,��A{x%\~��oc�q����}\+��\whI𗈃��Q9�@����g4ID?4��KG��QD��,��G��F������%9�G�xe��m���ȴ�B�#�w)�UR��GY����6g�<�j�n�`�ƸC����I��i��� `b���:���a�����F�>A'ӈZ]w�=^��#���Q��A㙟�q&Wf�-G�FE���E?����~C��gEj�,�l�v����ž؎l,:	pꝜ�Ƀ��*�jX8����ᅶJܸO*u4�ӴR>���/i-$xq���� �V�g��z̳H����Π��bG�8#~V+?A5G��O����h������tr�N�[��(׈��ӣ���+M��c�-����h����!���r��,��)�ܷo�c�������:��ۤA���A�L�G���W�񯽴���[B����L�M�e�ނU�zq,蕴�\b�s(���>��;Q^®Mf��itد�ڍ����k�Q�ns�Di`�%�ܝ�NJ��f�7����h����##p��(���;���z�����̆�ʏ��`x�+�<�I�A`ؓ��"����g�X�##��j�\���b(3��a��@�4ҁ�RW��T�xfW�kI��I*�P��R�s�t��)�,���VUP-�U�,ʔ��!Fƛ��^���a{$��@�R���eU��Z�X�/1*�G�>�B�|ck�2��������`pІcwz�Nt�2��G*J�p>�b�D�'�Q�u7f��܌��b~�,5DC����B�q�5�'!uT5����#b�
�u�{w�X\������x��(Z�މ��d����l�,3"~�����!�k��&�;�}*N�4�@�B7�A%�(��g4��\�8`G���X��N�������CM��,��V��Q~�r�Ο�nh	mu&;:��'Z���a���p�f��$��b,n����z�Eb����5ґ�j#[�iy�c@�/}������$��	��o}!�1d$�'aK��|͍.7b�Ž��6��qBt`��)}��Q����?~�F��1SǾ�����O1��!�:ֲP�Xm�����ܠ��+��l�0�GT�(bG����z�6���ޣh12�������0�:�8��CS�m߾��>�O9��bLr]�N4�}� |{�ޖF8��嬷S�r&���'����c�7�,'�i�/7�`�\yMb���L�RS9�K�̴��ϸ��3��M�ǵgS��#h�yDٷ�>�C9��ω�?&t��ux�Qg:�����	������ֲu�T���������ӏq�Ɣ���Sg8΂�&��X�vG�&��`p�Xd��"��v�s�.�|�z�2�,c!�ȐDс*��:R�r�s��ҖO��!`x; gV!��Ô묋_�'�@�7���1��&tp����G	��la
�ё9��q�!���*�>tVKY��F�u���)�a#G�u⠈�82�EN7���u���G8Q�B�,��a�K	��%����M����J�ӗN��E&�l�o�D�,NT���ox���ԥ �Dq-���#���潗�ǟ��=q�T�M�PnfM�%�+���������8�k{&��~�t�+0�n�� �p_�}��٧�S70u�|�q�ƾ	��x�[1��07�k�<�'$���6��JƤ�"���-g���r�	�!hM��N�h��Y1���(�C���KiF�D�\���
��H����؉�=IE�K���S~�L��q2�7�l���[�!����n2�
�N�-cȣP��Q�A������L�-@Z�z�9ʒ�ܸ���~���i� �?���c�6^j�P�J�¹h==�:y�8fo;�׺.��@�8ۥ�r��oH%��H���4��g4�T�-�S.؎� ۃ||8��㶶�����F7�~G`8K�"���1?s!�i�Ά\(4:������)u`�Ģ��g}���Z����N�L��种aw6`v���}�(���/���J7&�9a����ol�Q����7�U�1�����wsF�����0p��.ZDS�Я8X��VÁ�ttsP��~N�J3T��-I��Wǚ��/�ͯ^B�2�~��3��:%�_�Ո�����tL[ЏzsN �n���l�8̮�������\!�����qβJ� �+~���m�����z�/�&_c��Zo)�ؒ/�2J�{��atpb����k�p�Z��K01f^>�1�k��[:d=tA�w+�{�։�s�̵���V����`�<I��%��J=�h��ry>.�f �*P?ُ�b�t�WIW�}�W>�p00�3W~(��̵���j�}L'���m��n�1���Q��L�6�^ëwi��d墉��ĉ�π���|�r�c>���'����N�5S����M��l�������JG���Jt�ՙ��d��L��>iO�zv60R���8O:-%{�s��&����/��g>�M'S�##.Ap�:Ӂ���|R�E�<+#CgMu��)�H��(u��Ep�w���f�j���<���S>�G���&�8W��@#T�ƀT>A��˷�3h�.��'���!(H^`%}p�|����:�^܌_x�T��'{�5M���t���1OIz�S�-�͟��=q�d � �� 1`3�+nǿ�K�ŇM����I�QB6C
�ݝ��asK9�Ὗa�,��)7}�x��Fך������t����˧BѡRV��gJG�Vd�Ή�>�s��(�8�{q�>�S��
�P���=mʨ��Ћ�8�a���~k�%���k]�-'gk� �0\.n$!�{Ȅ�Ea��'�,�N]�.n�L˔��u#�?�LL��:���Q�>҄��
��SޣT����rCL�&:־Z-5��@4vc<�c1�E�ۼ��cإ�0�ͻ���]6?d:cň�	�	�.�*B?2�iM�T��5Ga��}�ҡo]k3pq���2��i��<�_a�6%�����_	��X;�7��\�w����KrI��')gw��O�A�
Ʌ�'���6�O]G�r�����Ekc-����V�wp�W�bx�����Oc����gq���y�\����%t�ޏ�#�68��(R�/m�K�u��#?H݀��hʔ�v`BIr�,�ANNp^��c��}�P���t�)r��2��
bSq���d)����*m�Ǆ�ӽ�?q/���f�k�4~�N��F����=�iupzp*ǧ��;pu�D?7���s��^j��u�A��I[�S��z/��/�tS#�0�� ���}9J�N��?m�/��D�٦"����R/��'�����Q����-�Z��ڛ��.����,�	.��`���t�	n�IV$��@�[g� "�6^zWj&!�`��9P�ܛj
o�p��#�5�tq�s���z���6�����x*J�tLIW~u\�e2ؚrŹ�S�{)[t��O�8\&�LP�h��˺rP		lw��"u6��<Pң��8N
��s S�r�<a+
/�|	�@���89s(�d������:��r�(� ���ˍ�n,�:������G�^��Hd�j�����:87�M?���o��c��~?��ǵ6�
줇��Ol���m(�
���:'�F�tz���r'��͍��k��!�p����������`����'��[��?k��D�,J�����e�ɣ��f�������;��~|��;q����,s�k��Q�.�������Qj��ɡ3R&��6�����數�(6g��m��Ο3,n6����~�l�DCa �3 �2�ܟ�bs�֗�z>�q֓o�pM&���שP(�f�WJ"�cS��i2nr$��7ft�H.h�0�Yu �@+�=�
�Gpp����q�td�F�O�L���^Q"��-V�!��d�nN�Y���Oqz�������S�X!�Jo��4^T��n����aG�)B�@vc��6��/a�0�G�?w6&��pm5b� �O��;FމuH�����~�U<|�Vc�:? ��v��H��F�\4<���nt�7z�X��r]b���7b�[���Q���vW�R#/��Y�Y�`ĸs&��1? /��������Nٟ��lq��,��jp(�VV�~�T���޽��uj-���G�O�{=e;�"�); o�l*��c&k�h��{~\o2#[F���p��8d�T��@GJ�rCTi�[_��8��s����m�ߏփ;��:#�?�z%F8}���^y��� �6�2�����:%���v�SG`�G>�L�������:��yse5G�$d�9��H�d���C��ރ�w�w��י"W\|.�pܡ�#���[��XɌ��c��t������]�@oaঃQ��	�ͳѸ@��B��v:Q�����/��V�>�O����O�Qy�~�#�y]i��C�D%��4q樲�7�J\n��u-�-�Z��$0�ZW�R(��CR�7q�$\�]���'�P���dPgs�aī�;�E\ꫬ,Cy)C'�8��@#>s�,�9�c���]�sD�Њ4���Rw	ݼ�½�3!�k8���%(o�N�|jc�:��&yM�ϵ8s�5���J=&�#��f�C�>�y��m�N�� � ͔5�$�2��P������u;��1�v��G�߬�N�">U�9�g` �6u��9�������~���D�S���Q_|����&���5E�_�!\q�vC�Vg?{�������6c�G�±-Ȁ��"$䋓	q�R&���?���nP�wBFD�����N�A�ۿ�a|�q�c%���8Љx5�ȼ`IM��I�%�	��W*����U�ac��o�!?U�h��]	�q2�@A�D���J�jJo�8�>�C�t�������#�\�#��ȍ��"�π��IZUnLH���8�0h �o�X���]œY�������C��ђ~ Y��3o����e8s�H�b
���$���4��8�_�L
���F~��v�E�k��n܈�N���X�9�YQ)N��F�Ԁ}K9����p,F+ 8�0�n��-�����(�@c}3&�]��2��~����n<�Q:�8Q*Ui6ְ�g7�i��a.���̫K1=�B;֣����(�{����Ǚ���~���l'��n��v4��'m��p�o���մ�'j���z��k<
�p]�7	h Od�>��r�3Fdt���!���ѥ����|�+�(�S�����Ƹ��|ߴ��
R�g3�.�hp��O�[�#Hin}�a~���_���)��M1��̑���ut��|
�s(�`�C�oEύU�-��ի1^�~2&yՆ�uC���L��+�zC�(KƋ��J��F$��A��&�Dso�4��M�o�f8�M�(wv��9�1��:����^�	N�3��{z8�)i�as�M�����Q,��h����f�0fØ��E����X[I���v|�&R鼈�Ͷu)��}A�M�P��|�l���@^���k��\�.2,}��� U'�ұ@Iyϸ�z3e�PN��U�9���m��d��qV]�nN?͏R'�f��3��umG�ӹ���l�Y��;t��/�8�2C�	��"O�5�SL�:�'�sf4�+	�!|Ζ��Ɲ��t��I(�?�<�9�4fP��jd-[.I����.��� ��q2A�O,'�	�{��B�f#�䦦�=c�ܺ�k�著�i�G��?�5K:x�*�'|L_lJ��������׉Z���G:�����X'���!!���<~�j#������ی�:�\�W�.f���z�W��D�~�>O�3�X�(C��wB���0"t�P��Wnƿ��[��.��n����x��}ʰ&C@`$�*���Y9v6�0΍����	G�6 \ɩQ��`1>�2�?ڋ����gw���"g/X�~��8��N��` �S|eW�Ϸ+r
ZC�RP��W�9-�H��1#8�(ېy���$䷽0��!��.�&#Ip�}��m ?}�ŴkJ,��S�(=ґ������q-�\��M��
?G�*/Bi��Z8�U����ۮ!4�Gn���{��,E�֎6�k`p�8�c��i,�#�փ�љj�`��a�u��ܓG\P�����WN��;zt�Zhk��F�[��ܹ�G�-?�G���Et��1�s��W�n�1kesE��%j���.rt��Ʃ�M@��h��h���������p�V�d���e�UHyy�]�ʰ�lo8ӣ��������j�_:�i�>x+n�y"Ag3�І1A*ǖ�+�5�IK*�Y?�T�NVe�9�]Ǉ`����ܱ8����Vˈ[G~����l.��::؆Vw��y'M��k1[ՉR?�O)}���GOؗR��G^��?��d���佔^�,�L��(�,���9��"�#�F:���Y��y�B���i����	LG��]��ۯ�G��,2�s�a4��<��>���y��M��@�8��)��%O{����m�"��pi =,R�%�ߝTݒ��ßg���:�s�ɖ�u��M�N�+���ȾH��}@СJw�E9�m曘��G\�BG7���P��;�,qe���r��W�fC�!����Ce����� �����Ϊ0ɛ��Sf{K~��J�/�"�I�:��l:��NMz���K��OU�:���/a��8��>���H~�.�5���$y��QInR��S����7ޜٱ/���g`�g��O�Y:*"���tZW��?�`Խ�|Tn[�>��������V�U��׹ �x�@<���-�Y���7��bw�Z3��7㧯�D�F�}�D�ꅯ��g��o�Kc�?ky�*�����D� ���#=�]���_�u狷����	'ѹDi����
!�(w2qEX;�:F3?��`�'X�^�@���<G��<��*�C�F�{XX>G�i(&1Ax��*3��Sr*T�MK��Q(��GG������1���?G���'/ ?A-?�+���pR8F~���N���>I���B�V�Cop��PN��B�\�+ѦuN�R��B�3yO}θ�š����XP�P��du�-)_`������?�:)Ԝ��>,y��ఖ���gH�g���S�]5@�
=m� ;O���~,�_��ga� ��>������J1��/�lW�rJ�����'�MS�P�6á�6����<>�މ�{�����c��rD���O�M��yfF���Ze�qu�&x���0��m���Kqл@�9ˁ2��LjGP�8O2�d���׉�N�
��tti��A�=<�ڹӱwٍ5Gѻ�$Z}�}��ՕܢC�����3*e�%�5U��'�#yn�K�z�:_y^����1����P�q��G$]}4;��C�NFQ� �:��0x�_{>fkk�D��=i��%��ȏ)��I�f>uPR�+�6*�f��F;@�3e��� <�H�������~������g?Lo�Ƌg���#�=<�_i�|��!g��F`�x�v���rpY�E��K�E�션�7��q��p�(�Ю
_Q*�ihH�l�2D�Eni��v���y��-W�))R(@��*5�?-q^P�vUY+Xyp����Յųzڄ^��*l3�E�,�'C�g7��Al�כK뱄3�l���v���dД�4�� ����W&������r���Z�5��	�U~Җ�5�z�]�f%r��J�	iKY�ә]g�ʽ:U� �"��nw����-U��$i�q�Z#7&mt;�d��4����J���K+�6q�@bx�5�	����.�="�h��[Y���� z�u����a��)7���-��oZ谥�n�;�vn<�&Q?}���m���؟�
��f�к���1�Fg6_$ �<'O����+�,@;��K�`�r�����6�Rw�x�������+�p��C? /� @gkM�'�����xZ��R����q�����e'��o�ǿ�����n���!�=�ɟ��<�v*�����h=�Af���ןg�h�e���V���Ly�L���  h9�P	P�����B $f��=�E��{����nG����aӈ�Sl�WE�|�,$#��X��ht|S�Z9���(}i�F�҉�I	��R׶�c���>FD�(�f��е�" W�v!����Y�Z��I<����^�xSyC�s��N[��R/��y\��D_�uR�
�;�����x����V존�L�i;���rjb�Uf�i���M��F���XE��(�i�|(7�+t�͝t��/+�}�KB��T>".gwP\4�{G�c`�/i��4��a���Z�/��ƕ�;�h����h_>MF��چp� J�7��F�s�2�@�}�t�}���/���(C}(F?�ܶ��Gb�q�,N9����6G��_.w�d�~���[��}�Qq��1GI��]�4N)Ε�LOu2a��UE���)�����տ[���4�[�(Y�rC�0v�M��W0:K� J�LwMC�3"���t�#���h=y�\�Պ�1][��k7諔_�Z�L({:��̍*a�)����u(��"�|:�ߌ�h����9:�ZG�׿�*���'O���I�醳3?0��g1Tϝ��`I�c�||0gU�+�}���#�=���#n?���$�o�~s�7N�����i�#eF$�~ ]8�����q�-g�3Z=$.%f���m)�g����ڄ�DU�H�D�淚+�%'�ˏg�?H�%<��	�&���KI�q���(^:Ո�K����C����S�$�3w��1���޴��~~um}5���Qҡ]���Gdn�7D�mz"Z�6���}�V�"L�U�I�4�{D�4{�t��S��	&���!N$�m���/uL�=��:���t0�ro5pw�'g����H���5���/�����i|�F�0��;:H*���s�q���Ct�<����I5e��s�iz�r�>�4���"�����_��=Ӈ���Q3>؞ģ>4�/�Ag��=���E����r�I�#��ױâ�rﬞ���Ci��~u�C��,/o!8x�x���?yy�Z�lA�d�V'�g��\'��G�������������z����w�x'n��'�ΏO��\�);�
�L�m�BF�dr����as�h�OR�a|�|7�F�_8�Wz5<�a5eb�6B�`Q��t<����J�k�0��ϑ9�+:9kˌ��&GG���`+�j́�~<YE��8y���mF]����W�i��ă�B���u�*��	���z0�Ʒ����t�����a`9�����&JI%�[5��."�D�ǡC�E����ȅ���$�Li%"(A�HC%v�������s; ڶ�ҋ��%�f|i������<gqdP��ط�|W�vw���fq��tƨӯ��*/:� \Z��^Nǫ���؇|b@��P9�N��W�QJsw)?z�q����;�R  @߿#.M�4e�_y.����5�3���&L�}�p�H�؏x��R�_�j��۟���J:Rl{��3z�uE)C����\"��t$\4�z��Q�<(#o���zvpp�cz�L�N�c�Y#N.�֪7��m�;n�bT���D˷�@^M �����mG{�Q�V�Zv��[��L��\����`[���ߜNP^r����.,x?V�_C�RVn<c���3)���6�_ں��>�9s��L>_�N77���J'�XY�d���@�����J�e�(��yssm���O�`��/\����}���-峞�|��_��Mt᱖/6���N����h���\�n�(,�aB6���?�Fv�odz����
�g���U'iR��E %o8[����RB��sq��Ć�:��Q����Or���X$hTu��m�7+-��zŭ^������ܩZt��1��͙j�>�7o�:3�B��#I~�ofN}Ċs\g��օaסq�+����'�Q�T���-*�|�Cyx�=�R=p�>u����r�*'�.G�IB:;��E�4]ĕ�R'Lҩ;��3�>m�x9�3�zY:�7��I���#�~�Z�����
x�~3����t+��(���m�	�N���yqu��d�r�Cx׭nƃ�	v�o�ĝ؈'g�D6��l�\�֫�J��&����ɶ����R�{y�a{�!��Μuq�~�J+���k�sW���Oq�hA��Oe|a��<�?V'
XP4���x�%�08�A�����ߧ�d8��o�� �.u�^u��2-y*�9eG؟D��X3i!�2]��ًM��'ί�_�\|�b˥#x�t#�U�arT1�!��T��j�!Q�\נ�`ݠZ���MI'q��I�� MR��44 ��Sm�yst� �U
�S�,N1AA􁑊���Tm0��ZVaZ��4��_c���(o�g�(�t��k�⿋4+�hi����!&"_��gn�F\���YX	���3��tM��G�0"k�R9�cy��֖��nĹ�?F'��[O�OVb�>|�>��l�Gȵ���#hD��k���n%����K������Ҋ�庆�F������J��hl�Ǩ>�5��>s6���t\�ޏ���"F������p�t��*>��F���}3�(��o������!&g�E����^;`	�8������-(FM�����:������#F�q��p�p�Z8��L��kp��(3��;�2����w?��/��ܩ8B��i�F}���D}��}����o��t���0���LL.���H���T� N:�K�r�Hoa~�M躊AuO�����c�������������㬔u��x@\�(U�X�S	9������D�}�>��7k C�ȧ=���D��n�	6\��O��׍ѫ/���Y�e����d��X'��!��-qE_LZ����Ѹ�8��Gc��6�q^[g���
�iѯ��Ƥ���"�PW��9�Ͳ��S�?N$D�l:6��E���9N�!g�� ���Y^�H�O��t��n&��ڍ�[P� �6ǳXe�r��j��k��疎�{�T:{�����wθe݂��m�q^@��ՙ ~�[�T�ǅ���b���&D�g?�&��}YȲ�
V֥�✚q;��E*�� �/��������mM]��1��Η:Ձ��@]��v�+0��]jz�N}3�\Za���@C��__�1�ĵ����� �r{Թ�@g��b�`�p\�[õ��^/��a'V;io�u�Ң��`�}'��|4+b�/l�@^6�p_�`@|-��"z�/6�_~%�8Xg�6%NB'�
lcw�<:Q���"��+Y.ٮ�Q9*��p�����8~����B4�A��Rz�)��{��#�u���5T��k��5W�z4��Q��� �pn9~�����Kqv��%F'=<yFm������]�Xm��\�����ǈ���T��E�^|$����
5ՙ��U8B�G�εp�����h�I��2o>�_�s�O��o��nZG%�р[^mO���KY���k�I�)��tA<?o3A���)gD>��w��a��� 'k��c�G9��x�1�}<ɼf�f����q�;p&����C���=���8����ܩ�h���;�8���砝X�͗3��55?�ځ���ȏ��c��ݨ)�^{����4�y�{y��v�qj������~9^|�b�z�t���18`�Cp�T46�q�@�����n(H{rsB��t�y�Zsh��O����-�Z-Gs��~~2C�3?���M�t�4.�.��qԁ��z�FC?t����nU���j ���l:�ȓu5@:�Du$]ӑ�r��}�tH��O�AS��|xP�}Q��_��:��L�Ӏ�<��!~���&����8�xۄ���zy� mrƂV����t�S�L�����uguB�f���+�I<]0<E�h>ي�ӧ1�j`��0���S�����"�@�-�<xa��������A��o�oϗH��1�����-8��|��ѩ����L��j�*��XD~,,�@��W���,�%qL�^���l̉PEi��ڼ��85�ʣ.N�U[ ������Dx�6�������ď�7bsw7����G|�ܬUC�@�J_��U娮�匆��Ш��>�{6��J�,��4ꜹќ�!��Ҧd�r_�ɿ0��q����צe���PI���\8�NJ�I���Rd9Ҏ��P��<���������?qP����J�S�S/3�#��s`\d �s9���嵗�7��˯ut��K�8��ƈ;��x2nc_�A����9'$$���v������R�$�_ڟ���V-^`���F;^��Fǲԡ<X,�,S�,�?��m&j
8;��6vP�0�$��݃�w�x7n�K�w�W�]wM�K��FjbR�<G�r��9���ߠ��1��G��-������|�t���͸����^*���p��0m΢`̊����BI0P�329��C��0>�T�h;LOƲ=�Vg�P���E�]5$6��Rj�t��|���P#�A��wq(�����U`�O�!g��ͼn۩Qu�kZ��#(�}�p4qF�k�Nm�@9=��0����sg��I���#>�ܹ�<^�q>.}����s�����q�Ɗ�M2��i�N��I�\$��I_�'�,ꨈ����3PIpRK9�q�Ή�A�������o����G�s�L��{���?����l�'/\��: ��&`.�Nc��c��](�87q�k�9Nd?�<<���ڏ�?��o����������Kp}	��B�����*[`���lB�C�ԓ'U6������X��~t�w�ى��^4v���xm��(wy
%?Fl{w8w0v��o��pb�N��>��gb�S�u��zO;��Q��=���^Lר������_��і霶��v���b�pTfwn��}��� �{��r�x�6����:a��+O���l����,��T*�*����F���.�:J�V�z*2���'�y��k@Ɲf��q12��1[߄J+�G0�4C���?r �fܼ9&N��(������$�@3T�^��E�Y�/�o��H.�<�Ub�m9n�"P&�sx-/�G��*e�ԗ��d���ZB��ěo1��l7�������C��C��ns��=}����R-��/Ǐ^Z�k[���G���=�mt=i�w�=��z��=n�%G�0{�}��l	�Iʐ!�g?�gy+툙��9�W��U����t�H�_�+Z��Uc@B�,�||���^5ﱾ�R��㝏���e(i;п�n化z�F�A;q�2x�8[��(e!Ar?s)Dw9�8,5�q��Ӈq0����f����;���p��/�� ��8�")�d(�� ��=��K�����$�E����k-��F�k��L�IShU�&�*̫?��m&��cı�w�k�?8�z;��k2�\^ҡy!Xt%wpnvpF�q��YG-!ڇ�\����_}q=n��Ʋ��_��r��=���ɼY\�72��>����$T�R�8갑�F\0]��Hσ{?C#ӻ;�鮧�����Z(q��뛊���R9\�U�4y<�!@Yc�N�|���Nm{v1p��� �7�4�\��ƻa�7?���m����y�0��u�a�r�K�n��s�һĻ�����첋@%����v��\���>��3�G�.2�zR�~�I�u���I��G*>������aV�:�6/�V�6Fw�V�v��>��ԧ��鳱���ތ���tf+=�0�Ñny�|L0�I<t3E�(��ЫI�\�T�"�Mڸy3�]�L<�ߊ�޻O:�jt�%��j���F�Z��e[K�mη �8�*����Ol�s�K���e?m�������t��=m���us#XF�����<��=�@;�]x�4qh�i��S��v4����h-Qf	�w��V�]�М6��m�י�	���6wp�>�Ɖ9:���N�����M�cT�H�ǆʮ�ۖ���N�#Ǳcl>2�6ohF��^F����)FB�"��v�����G�¹��W���ݱY��L�ܭ��y����#�ǌ����[|��/������ts�,.�lZ6�؀Z�Nș�r���	'˥��z�.Ҏ�;Q�q�߄eH�d>B)]e�nr�B�E	��������x�?yc9��1���|�K(�e:PǏ�;��o`�л���Qt��:�K][��3=�u�P���ǍΚz��q�E���N)g�,�^Tߚ��Cg~��:�%	��y���[��[ع�IG=�=ƙL�^�~��mt���Og̈́���YO[���d����/��o�۹<�:D>��tF���iO�G�m}8L�ؚk�࿚��-�����і�n�H�эo���(�Pp~?�H�ȥ������.�#����*�t*q�����H3p�xa�����LT[�ή��(����}������UFN^����`w�zg?v@ܿ�Q[+�0��M_ܧ\�#H���s�"��D�cy6�����Z�e�Xc:ր��)��+8%��|�/<+�#��<�,s,�3��+���)��1c**�ZjG΅�̧P���P�,1��r�O�r�8����~q.N�i��9�8,��1�g���T�!<�n��q:��2�:���_�U	�:+�-�	[��yY:u.n�g��'�g��O^�:ɑ�]5��l!�e�\�]���?3ZNG;묔����7���C�\��]�QH����ߊ��
�7ע�����\iϫ||�k��|� ����q=j�������7���h����^�(�k�M�G�m�q� q �'½_2Ї�X�'i�����<�ArQQ�|l�ԍ�z7f�\��},�����ux7�t���r+���Uў�G�>j�M'1����8�2�lY�½�湅���C�c1����?��e���ǁ~�FrQ�u���8īr$�lw�g�����I�#_���L�B.��4�O�Ҙ͖�H�8�ӳ�#pz�M?l1�Y�^H�y,u|�!�����D�!�s�OÏ�Z��ճ�Kʬ�XڀT/���`�bVȐ��CA%�� Lｬ�3T�-ҍ��G>�Ϭ%��*���,�ύfх�_=׉�܉3M�C�έq���;D7�)���:-�M���c4�Э:{P�ٵgx<ﳌq�nщ�>uz��
C$��1�ɲ�tp2���GxƑ�L�-�\IO�h�r�:X�Ӂ�,>EoR?pz;a�_�y�*�^a!/�����җ{�{�@��Y���p|��8q�AG*�ܧc��	Ǫj��U�����(�B���Є�I�蠔|��d��������{�wMm��]ބ/mO��Z����z�D1� v)`~�V�}?���!�Ą� ?�Ӊڋ��J4UGEC>9{�{o�͑���;�X�3{e�����3ז�Ǯ����rL��9� ��B��:��aQ����$G�Xp��"�sa���-�]�V�d�J�S𼯄��S	q��:+�D<�0ba�#�
��G9��e�p<J�y�'GDU��!�q�P@����p�\W�T��rV8��H����:K����7aʬT'g�|��ZZ���r,�H꽥�=�ƽ�V�&�B�Y��O��=����D�E%�m�&�X@�����6*s{��Պz�����:���=�v�w�PGb�QN��P��tz���儣Ñ��hW�7h0�� ��f�]���f���V|��{�d�A���Ά�d9�~���t��yv�C'��4�Q����g�}_�'Oc2��x�>����e�u�uv���_����{%5>���<e殑�����FM?6Kۆ��C֏��4l%?�qe~�Fx)3�e����ى�ߌ����h2�i��3N��� _v�|�^�`wy@�B�Q�P���t�0Mg�}/p�X�����Iq�p]��0�ݥ�_���T>z���1q��\/d�A�G��Ҩ@�\ﴽ���+�RR���FL�]�)j���M�ȗ�)8�*�ң4��L�؞���;.	&mJ��7s[�G_JIÓ��gHy���Hn'���ߠ����*wܔ���ƒ�\����4�N���vl�w:]B~;�uVĭDjNsB��sP�<�H�(4x�{�����ɀ��%�6�y���G�g~��Z'go�[�}��Uu��#R���Mڢ\�Ñ3C�WՑy,��>q��/ʧ^�.eН��繮#U�R��8�S]��G��R�<�M������8JY72�L�� ���)�+9a��ҁ�m�T�E�� ����6� G*��qVѾ���UƗ�����I�$�i�=�k:�,�D]]��+8Q/o�끭a�R�?�<��<��;Q�)K�/I�������❃����Exv���(�^Ě���;ʙ����F�q�6��~n9>{�Ln���G4��4�	
���'�k�zSU�#��o�r��B �͈K��qd�לS�hS:F'��y��0�{����*�ώ�b���2�Q03��9�(�R6�&�g�:J��Y��>��,W��<)��a)����%>�������z:J�O�J�Ƀ��g��;8#K뱊�5�1�`�w�����YT�JWz��n��8�������2�.ˎ)�:%M�x�]Bc�^�Xn��D].&(�	N��ћ�ع�q�����$�F��Gu�F�q:8r�Y����-��Q:�;˱;���p7޼�4��X��xٚ)H$�ն,䀓�:��.��yַ[>��Qq�A�H�+��(j������v�v�`�zLz+�����qj��
 |;Ĺ�����b���8C�w�~28l��Y̆����Rԇ���r'?p;����i�ܔ˵Q��|9��%�iڎ����~���2�\�.�R��ǣ�ѧk>:��A	K����+��AaIT��Ί����pq��8l����qݘ^���g"��}3��l��ц�~Ƿyk~o�MA}� %2��$��FdV�Wb�����skѿx��Y�т�j����8�A:H��_�ꁼSg|��B�Szo���S��x�,�98�|�fR�)��8`T��Qr���4Y�vX�7�lΦ˶����p������Ed�ފ���M��q�iwj^өArrp��Q�[�ʅ���0u�g�i:��JO��E!m��Z]����a�y68Ew%<`Ug��Y�\�`�K�#�V��e�'�*�T��J=�Y�2�V������/�՟::O9�.p��ҦR�NQ�7�:t�r`��E��-p��O	t��K���dvo=ډwwg�3[�)z�mZԒ2��Leٞ�u蓃��̓|����.L��@װ�t�V[��F7^őb|w̧�+LXy��?��cŠ��ճ;w�]�5������N�:+��]�(��2*���D�.�.�K3ZM�����q\h�:_�2�n��z����OFᨪ f�t����x��E��_��ҏGZ:5���8�2���1�T_���U�t�����<!T��P�����&�C!�>�w�<�W!���ə%���8�T�6�3�Qh����Tq͡��x-�"�9;��Ǳ�S�gy�sSI�2�_��=?��*uN�N:SƖ���S�G
-����FS�g���X�\���	;iچ-}�.���5�ȏds��\�½j #8���s' ��C�>�m��7�r���R���^ <�Դ93E���uh�M�^�) /�:RDO���S1_;K�N��߇$���0g��e�nR: Gj����gp�Č�9��؃~:F�`�d:�����y:DgN�t�bܟ�W*N��Q�wvb>�I�n�;7Τ�9��	�-���ߩ�~��F������f���q��]B@�nZvW����u��?����o�}�3T5_��t���h��wg���}�g�7�B_�YJ��Ǔwh����O�݋!u��x��uw}v	:���D'�z��?S��r,�BWy����-�y���V�Y|�#��HϢ�籸�������{o8��`�yHԨf.w�H���o���o����#"_$ ��¾Щ�ԃ�!���o^�=�NE�>�.����W��y�|������Ѩtk�YG:���@�9@Z��r�ϼ��rTuP�� ���m\���	��G��t���٤�Jǧ^s�+�%���}3�Qqo��L��`����?:M��c���*�M_֑m�.iK�T�l@���Dv]&J�P ����8�3�J�>
"3Qv�ɳd+��X?��� C��w�b�o��R�W��S��4��J�������'X�zT���D���7��g�n�golbԉŘ��>��h*U�ˀ�c|�C�Ź�jC��2�KRb�qP֣D�_
e�"p&�<>�T*
���[pТ$���3`UzIUu���s�w\Nî���O�"A�d0ZM"r�C�L�P>*TAz�8���!#=GO�J#�S�q�h[G%��T�O���n�8]��0ζ��U?_�oģ���]BƊ���ҏ^H��[	��F򙇾-N��#�d�����Y��A����y��Ͼr9._{��Ѿ�ѷ��u�ӳ��S��\fd���X��>͵N47{4~@!�m����Ѱ���X:󩸻3�������F��#8��(0�*�?$O��� �j{)�m�1��)F��19��h��S7��������V�5G�����=�:1C�����]��C�)1���^�r
~N��ޓ�-���j�"�f'Z{[ў�|6&�<��'����kC�#؆���sc�u�kN��A�kDk�����vk8>�=�<�sm_�@�}�����5w<���)�స�Ny�/jv�P���Go���~�Q�oC�=�x�8z��w�}��� g���H�_n����mGs�^4��Ob�����c͆++qx�<�8q�Ws�#-9��+����҉N5���>¿Uȸ*{������/}�<���cޏ�V� �w�b���0�,��.?�g=x�NY��v���r=>um3έ␏�̗|H�1�n8��(���:�ĥ~�z2Oum�H��s�u��z6��(:2����Uz�<��Rg�V�N�9+��*��G!�]R�
���1��re���g�iy���2�̓iE��{���E��x	/�<8 E��|;S>��X^���y���ͣI|��n|eG��hL��  ����4N6�qP߾�\Z�љ�����4Hg����v|r���3X�F�4K���G``�����OT��D�"HG�<������{�Qe*���
r��|�Q�<���QV���?�1%<0��� :��qi5���R�8�ø�c�N(�(��������+�@��d8����'��\���δ�`�3���W��BF���msi�?��U�3��U��)�D�Y��z/I<�kF���<Y�R��lr͎���/9;b<pk)��!�̅�������.u&�M	��q���3yl�lp�5���������$� G�E���<�W@�}g��B�����^|Ac>��M��(6o}#~jc���G����q�:1=����gQ���ҥ��p&ߌM��$�/�����=��3�a�q�?i���˱|�����7�?�o�����E��X*?�L=��� ̑��,�x�<����	u���X���G��H6�]}����$��R;��=�ӏ��s1��C1%�ux'z�w"�c䠼��9�m��b�4f�Dg���?��7���;��}��4�.�cs�0�č���;kl���gb��D��עy��R[�����\��U�Ѭ��[F4֣�S193ꇷ���N0�kv�r�0�:�w���љ�1[{)�F�<�J���ͨo=ŉD���i�Щ9C"��:��`��]�4�G�ίGk�K~�ӣ�n�����#��g.���˱�܏ļs
��Q�����k,Aq��]1$(t�I�:�q!��r��'���/�ɩ��|�{���b]v4!eUٕ�<�S�t��Cnq�1\��".)Oɢ��F����i{7^_����^���q*fۇ�=��_ɻ�Q(\gW�휙uTm0$�@�)�^I�B	���{i�`2M���
��@� U,ܔ�)���L{g(���dX�t2�����Ԗսyg�_t���_��:��tC�,����n�����QK������v$�ĭ�6b9|����?���⋻��/Gk��!o���v�*�n��k?���6��d� y���f2z���.u�__�_��k�b��0�W���ߓ��:*��L���2><�Ư�AЎH =�S8{�U�:M�g�R`JG1�i���\Z>��ʸ����7�U�O�	G�jTn�
Lx	>N�H��.�8#���Q�Z��ř�BN}29���䈪�s��֞L����P�-�E��%����k�Y>��+��YxM�����E��s���Qe�;���§�#���׎��Ag�,�x���d�"����q�wߡ�S��N�Ǹ9���B�)�ҋ$���TXi_���2�l��ِ9i�JHW[�nG{�A��4�/�v#�<w-G���AL�|9�ߣ8����h\Y��<ɻ�UsW���r���#nE�C�(F}|���h�z!�|�n|��cۭh;πG��IT��Ĕ{"�r��Ù�T{Oދ68��>����h<����h=��p;�㭨=���Sl������}�f�~;껏���0��be���N��\�p��ߋY�m�D�ћѽ�k�޹���ўn��l��i�w��mEg���8��  ��ߊΣw���q�4b� �#`�mS�tڍ����}�\�ͭoG���DG�����Q\޿��y�w��=�o���t˗���Y��j,=�V�����A�ԏpt�uS7mi���Nt�К��nD�6�����>|;�{���ю�h�g����p��1�^���5�����U88["r��0qɳ�'�73�P����d8��rW�z�S��_jI�_�[\��w9�sH�ޏ��{`3O��6�q ��mst�O�Ĺ�&i.q��b܄X&h�M��n�:��:��3����y�^�G�]�}���R�1֤��8�g2�Y9K=f2���.y�2*�s�f����Gµɂ�����'�m^��&s.m/��3#�?g���袜��X�����.��p�.�~��n�7�m�c���L�}C7CG1�T�"�;�IF�6o��E�@_�:�A}�Xk�K�h��I��v�}����I��['���$���׈��0/�.�w!���NX�/���e`�YG�G���!������܍��dY�*\#��Nf�z�;�&��z��^s�<�s:c0c08��u�3E�LC���q��F:��X^���N������)%��'K'
z�qQ�qe�u 5�ɔu���̗��u���I�Ce]@\8O��r.\7_:(��J�M>��+���s���uPWV�8��o>��߻ݏ�C������0����c;�-ఠ�I���"�@=Gs\� �.���_M�Dg�v�l�g^<p����t����r�\[[v
#�,��0���.�d-�q�<�1$�������D{��8���7�y7�x����� 9h%�
S%#q�*�3��3g�����1q�n��0N�w�{�-���G�'�#����Kǔ���A���F��X��	�I��G�8	G�I�JtmQ�>f�3����G����q&�K���|k�(�{�1�>�����h�o��8S�����8?}5�	�4jRO}����4���� ��:���ܖ��`�h;j��}��q�u�ɧs���}��7|��o��F?V�����u��׷�\��|�	e}�� ����ݍ�kA�g��s&j��o,�~��E;�8����s�\�M�%�㺱tn�3�S�|��Ic�_B�w�(a����S���8:�@�Q��E����c���w9���e��7U��?�}Q�A������ӣA�ot�t������O�Z���+J�`+�B�h��r�A�H;���6�/⤃:gq��j �Q�w0x��$��s\�וsB�e�K����p>qx�#O��s��{g:.G������n΋5\:Ky�s��]ך��BG�>Sz�`8�5�����pv4�߹���7�W����F�r��f�Ͼ-��0wB�*�9敌J���%�C�׉j��:����f���$��f�����}�7����~�C�"�Z��Ŀ���'��%����2��!�+!�&�� ��$�j���o���R�u0c$y}����F+�揿?�k(�vN��)�[�~p��rEgg��%���*D�׉2�(�V�N�"�'8OH��;n/�[���ɐ�i��]$dY�Yݕ#�&��]��B�!�
�F<�Ī@�@?�.�#�ė_�|E�%)��9���`�s��ةS�đ��7���\�f{x4��?؍�������n�����	:�JҧvG�ɵN/��v���Dy	��npk�j=������xy����WO�>yG���ˣ�ǹ�-�z+�Y]¯� �Lq��J�Pv2-/w�Q=��Z�xr:�?잉���7���Ɠ�i�{�6
J�|����f�-�/|^�s�W����0^Xřy�7c����r�	N�o��5��Tٶp\W��q� Vqd�l�������1����ݏk�짍�����4�;���݋�gN������~�lu�I�EI�;�ku���9�`�p�2��;�?�Χ+�� ���x��K�t�t��h�0���ӱ�㺵�8��|�qv?*�2���t�N�/w��^8���S��m3�|����8i�Vt��0ƃAЍ	�?�^|��t8?��}h7N��w�\�M�N�*Nt�Z����cp��v9���38��|��p�+ e���������ѕ>�[�2i\�P&{ݜ��U�,��l�q!q^g��DVN�1l�����J��+�ĕ2:(�>8�Iݍ�f����ꐷ?��� ��'�����_�O�Y����=J�� �2�S���-Ucu�8�ձ �٦�T��`��U�7)��yz�3��/��:/�qR��>�ՐQ�X��`�q�S����ź�����q�%#��#]���m�@rH�t�ISN�������|���+��b{�,��2B�fDg���eY=p]�)��Ǫ��Z��O��ȵkn���C)��Y���z��kK�\߈���Q�����>Э(��>|��(���ې�NԿ�%�(�D�:Wt=�=��
�|��8J�,Ͻ��o�al�K��u��qv�I��O�����ǋ6c孑�R��Z��,��� uX2qVX�u�L]gn����ʻpS�3a�`��xӝ���𩄉.B�����B���"�g�@#i�!���l��c/�d�?d.	���������x5Ig�7Il������q�_�5R�,MRY't�ȫm��!��ً_��_�����Q�Ͳ�(Zc��v���BHB��ʁ�+���o�ə2���.`v���7q6�t���;�b��o�s�'q���g ���-FQ;�h��+�;�f����Q���;q/գ?Z��;��p7���u�ĵxrt�8�5�(��H�G{��5d8��n1�����G�g� �� 6;�����۱��q��k��k��י�e�@ұ�{c]w���p�A���ĩ�p���i�9'Ɛ�����P�ǣ�Y���wcp�4�^{!N����<���6NI-�k�i��8����&G{�N���f\{����o}=��u�����L �8�^Z!�����xo/�_�+��ƽGw��pZٗ�\�q(�:#���`�)�8�����ʥ�薈7��v,��l��������铧�6���Q?�{[���/��6���70�X[[�8]�C�t8pvG���l^�����>�Y^�!p�2��.4�>u�a
��t��<�'�K$�|3
>�YFY_��F�
�9^���YLc��9Kß`��:�1޲UT	J�|�ѐ�R�Q�^3���5_�p��C9�މ��ø�:��^��p�b\Y�D�^괔e��g��$~��ʗ.J^{�h��	����.3.�Pp-?Y�1��U�vA�&>�/2|�X)t@�D����NT���'y��2�}߲�2���lW����
}tH8�o~�4���~���}Rk�|]��9�ʯtJ�Kx-�;@u���.io��p୳�����
 :Q�Y���F�+7z�^A�t��w��ԉ�>�>�3'j��\s;����� ��/=�o?f��t��pd?�QJJ�y�7��0--��à��qt'�8n0��R����ӧq��Q����������q�
����f.J�7�r���=��c �"�S����&zQ�Wޘ�I��8Z3rq�D�7y�U��wa,��l��2���K�t-M���<�U*NUW9K�~�$O�/�ԝ�djVw�]rEX�Dd�������q���`�����̟�yGe���������[�ˏF�F�__����1q���HXK�.�Q֑����T7'C�G�*ib��O���ȭ�	��I���v�q0�Y̻�0��؍�l��'�o��}"m�ę6qXs�F_��SOHő�^M[q0Fn�X�:<��~�<xLPKg�Z�	Q�EX����s��P�z-� �Ԟ�s듸�Q�������_ЧmgNo�/\���w�y7<x����8.1��v,�����ql����ʍ���+/�'�o�w�?�?[�kv�p�AGq��X]�nߍ���q�W�v㭷ߏ�?�0�r���ǉnt���g/_�>��[�މ��V\�p>�\�#2���q���t�|Sj48����磳��ݏ1N���Z�������?����m�d����܏��]��\\�|5�{�gOoĕ+��O��k��7���A�2�f���c����ߏ���&�Y���)�
��:�mӾc_��n�S��v5�W>��}=��r�O��5(8����:��y�V��ce`�`�k�Tf��e�(�U�Av/N�R���O�U2�~,�C�	׳����?D��-����2���uBʗN"$��6v�Ƶn����ӽxi�k~ʏ��ѵ�Uǎp�ՙ�m�Ne�P�(ۡLkA��8�<l~�2�oݐ2K��2��7�]<��p���V!��$�Ҝ�'rX�1�xN�\��i��z�t&�6�B/a��0��[���ʯ!�:��Y�ȿ lc^$��,-��<���yD������(�l���Ǘ�8PK1��+��h�1d*�-�(%������ u�8C��3��~{f��eR'�eug��FW���v:Q'j�(u9��
�?��O܉2����I@���gOF����V����@'�ƨz��ډ#��7.�Cy;N98~�e�&`aSG2~>qOFjxO��i�����9؉��8�-���j�r��#�儉#�ѝ�][��Q�V��y$�S�����D����2����4�|��!�Q��L����SP�g��C��Xm[�k�ϏQ�aV�aD��*d V:>��^����W$C���U�|�&_��C��G�8g�u l��	��X @�/�(�w��h�M=#�����0����!�̚�  (
���DAWh���}�i�XW!3�㪒�\f����Ik��-|���>i���Ø�J=���(�x���v5Ex��}6V��z������MFr�}�!�^I�*�ĉ2�r6�x��)��pԫ��xp��??���b�7���ŐQ�����7���˱��o��^|x�a�����"*�}��^w)���b8t��N�.�ⳟ�D�|���F񵯿��pG�NO�4��S�cee%���Տ��+���_������_�ҧ:Q�XX�mnl(��?��p��B�:�������߃w�[��1R��c��^/����Eq���x��[�����7��Mp:
_��Dm=�κ._�B�K�a�x�����s�8z�Ν��y㝸�Ctϙ(t�8��G�kƥK���w��M_�r1~��奕x��o�w+o��<�;|7_����ϣ3Z1���8��q���p.�|�]�n㌡Q�K�goG$o2�K9�.k�<o�$���h��5<�#�'4<�cTr��J,��Y�+�oi�(]��/��>c5�����b�ʜ�mvi��#�x� H�^��"pRx��-0�|dR�HS�t2(����Ò.�~��[�+�˙�tr��AH�J���K�1HUWu)����}�� �t��.�8PЪ����`���v���Ro�dӒ7tJ��3=�|KSVⰀF�t�����\A�[�f�ː~��A�O��џ�b��#�}�/8���_r����Z{b���#gڙ���g��ct������F�v-~�r/�ڍ���]^�U_�\#m��t���'*��'��$?|ik���ڊ��`������r?��A4F�hϖ���.z���[�ah_��?����	�ҷ�`��>�Su8d�1�`���Q�#�o%��MJ�L�_��1��.��A�-2O��e�����X<�9�E�s�V�Q�̈�$����aT򵺴#���:�6X�Ô�:
�yL�l�:��J=��/�h�*�"dv���f�UѮ�o���r��(��e��%=�6
M1��q�h�UtֱÝh��~��=�1E:�0�
:?ܩ,��,�X蘣7�$��	��rн�s�bp�u��t�����G�'�kifC�����Ǚ<��{�-���������Pn���o1c\T�d�OG[�Q�@ׄB,�]��Й�-��M��/�������׾����O���LF���q����6���[��w������AΐJ���kw�w��1�����ܧ^�N�[8UO������6���n:[.H�vbye�e@ߌ�'�3q���7��0�x�8���q���ۘv�,/��E�^��\\�|>�v���Gq��ӧ{�g]������E�ۦ�.8�cmm��<��ӈ�G8R8"�̳��>Y��p�|��p�[��x�h���a��������9�!��.���ߧ}����Hgg����Ƶ���|2����h{?�=x�`�)7�]�ѹ����l#|�� ������u?��G_�>)h�|�|� �{�$-�]S�*��s�!͔<\n��
��a¢�N������7a#�ג//�RQ8��xp�F��9�,e�k?l;��!8b`<6M�s�V^G>ɛN��H�:!�,�0|��quU���k:5�(��Y��o���/���G 9<������T_V Y�e	��Չ8��ڛ�����󧎦��4��j�x�*�%�ۣ�HZM��k���h�O��mU�D9ϖ�%.^rC0��w�@���>�� ����Pm���W8�9x�x1��mi�)�G�CA�|�TG����.ǿ��r��n,C�-4��3J}��5V�!{]G�����4��>��5����3�PLܐQ��gѹ�s�/㈪qv��9
�/[ \R�R .��_�ύ�0�y'�kK1�(�8R�Cl#��3�0�2�\��������3���ev��T&�dB�e���X�lYy��!�H�qJ8a�HD��ų��������P寲���H'�8��*�|Y�s¯��
RR�:��I'�(,�}:%dr߭��Gͅ���D��[���P���B/[�#�Ϭ����8����P�s֛�g�&<[n�FM�o9��dF��'9�W`J�N�����m�q*�>v��'?���O����f�\��9r&��Nھ*/��αy��:�n8)��}�éҹr�B����������������k�����8���n�v�r���o��/��������Gq���\�ę�	�Mn��|;����?�c�߹{/�����������R�P���j8U+1��78Q�����g>�����׾���ߎ�O��_�ﵛ����h�ϙ/	�釿�����?���8~��_�Iē�{1��--Y� ���S^ܔպϟ=��̫�����>���a<x�4>~�N`q�v�����Fl�od�oo=���'�������j�����)Lԉ;��Į����`?�.N��e:�8���̧������o;�?z��֏w?��%-G�1����=�*�zLT�[���~:ٖ����7�µb���%g�.��b4��#Ne���t�ɇ�P��?|P�r&
8ΰ'�+�	ULK�4��}	՝��Z�t+L$��u�kv&�5�����;�Cǜ)�OZpX�v��`��`�u9PTo_��
�ͱ|�Ľq6R���ŏ�a�~���'����v��t�8*��v�?��r)�f��K�n~�W�th(���ڒ��ȳ�-���ʑv&�:�/�����f���_��9�Yt�%�,l���P�v��?x��N�}����"�J� w�
>�-��4U��>(8f[��D��Ϡ ι1�ycg6�񯿸�r7>��봇��d��	���G�}��;ώ����1�z��ϵ_�ס*|o'j�d.��c�{p]6�,�)dW���^��dL�_��&1n�a�!�f(�^,�W��\���V���o�t�ڻ���׌,��S(>)�5�>�"ͯg��Y�˫���3�A����-F�~S��.yHk2Rh������ �8��+������[xP,�|,�9���4p1ޏU���2_hc�fZ��ܠ-��m����/es�kݖ�V`ZƼ����3���p�ۇI-���Ki��(>29*M�'�������6.tN�d.�?��(��a�b�TN(0�0p($<2�^�Ylp)��g}�8xM(k"�?�:r�Og�O��W(�|m��s�f#��M]��.f��=C������>�Rޝғ�P�֝�xcxn^</?w>��{�k�������ĩ͵�+?�����~*^|�f�;Gb7�ܹ'�lf�9s�-ʺgN��_�ٟ����瞻D����o�N���XL('�8�Q�.��+����/�͛/�@'�������t�o�1em�Ϋr��O�?��?����qv����{���F�A���$�Fh����s�~5����L�|��X[]ǉz�>���7�Gg�4�G}g�ƴcϞ���x�����rm�T<|�8?~��K'�m�H>�����+/����_��7T��������в�t&j����9�}�:YY�-�����y򞏟�Oe����֝�d��'��o�X����?r,�x��x~�a��K�l��JJZ��C�����JY�6[F�bY�[��k���:��`~p)�I+�������(ч~X�đF��:�����y��\� p����4���#?V���ŉs�$�{�N\�L��6?��}u���,��<a�g�A��8��no�u;�v)�M�]�GD�z}��,�j�qk����#g¢v�i��L��oLIW���_M��luv\N�K��*���)8�M�Γ]��o.���g�G����\�[4O�O�"{�Oo}�뙂��7��� ʅ��6����6��W�u�G7"V<盪������G��ߓ�7HRv�|�����҈�:��i���C%��Ne\z���D�s�������:%.­�to�V�.m0����g$P��RMQ��I��1�X�O�~�P�..��母9{M|^O�o�Y���-�����{�L���N�������#욟�pQ2�3p��M7h��S��"���@9���@ٗ�8�/�@�<U>�#���i�\1���q(!��əvG
�g	%�_��ig��Y�I�<{/�>�rA7#RgU�t�7PA����<v�h�(��k�s�5�'�Q�m1.Gt��H�\]��\2���(�juL|�B3sb�WI��Q,l@T.*Ŝ���L_��� ���n#���ϝxp����=���J�<�q\���Cl*�*/��ɪΎ��J^�����Q����u\����^�|�f�ȱ��k�(��(�|�Ʈ�*��&P�����������.�	�ܤ�-�� ^!+R�Q���7N��cy�v��C��-��ԁ��<*OH�s�.�'?��x���4�}wJ�s�L���p8B��CwǕ˗�3��t���K���G�=y���^\���I��*8:<�����cח/^�Օ�lנzԘ�]���=����Qg�ݍ���ƕK�p�~jD����8s�JtV6�G�>��ei#�Z��zsH�JF=��`�4$ɠvȉ��A��T��Đ;��J<J�tpL�8N[�I�$��\\�DƉ��ȃ3=�gq�7�D��T���"�RRʖ��?��G��5����p"O4�,� �dr��-� u����r�1Á���䇣�C��{��L�V�2�0�m��i����KG%�s�s�=��W��N�~>a�1S?��&u$����a�;���	<��@"'
8\�8�_f�xu:�p(�#&���"�\4D�s?��z�<!7�ѝd;�k)���#����E��C��SF�OƇ�����{�ډz���&mh�ٹ�a��	�)���)�����_����]g�(y��Xk��8o�Y�b�Ѝx�7�U�0m1U�Vtu�~	�:�!;M%Bg)z����
n��?�YS��c���O�tGO��Tix�88�QY��/�r��ZQmG��
��5P����:L߀����}!�S$�|\TF�Ӣ�R���5��1DUFP��`��a�$�E���u���8��L�\pF��N�皉�u(;E�/:���A�|�`~pq����b�x ���y�NT<�4O��N+Xg�\��u"9E�pNp'�
���n:f������;hD{TF[Gغ3$�4`xH Y��}�6j�v�A�_ڤӕl�eHs�����3�~���;y�B�pq��]Ù3tЬ���i��{�w�/��	�N}�9|�m�M�6F���'�8��s���. Ӏ�0��Ќ4��`���~o.-s�b��	�oh�GE'�`g'�n��n���u`t|<+C�|RU�'E^�~sM����P�M��G9�p�
rX�I^������ em��8����e�۬IS�O�'�r�l+˫���	�cpx���'��r������z~Yr���2�g/��t5`C�_0�H>:��pV�N������Ay�V&�yul����c0#�:g���XZ[I��n%��՛Ѿ�r6�S�fZ^�5L��������1e��Gڝ�|��"�)����rNC��B�l��ԇ���E��K����C�W���rPN@��Z�����d��by�>g�8(Rd��(oB�|�;a��W��!?y����������5hS6�,|�r����{
���N[Ы�K|�8%�J�Y:8`+�0Ŗ�ef8����:y�r�����w~�R\iK�j�g��Ls��MKT�iȏ��rxj�� =�{�щ�D96�`�Rw�-�4Эy�c"�ӯ.ݕ�k��hK�n�W����u���6�:��+g�j�1���������\u��o #Ŵ�tp,N�$�p��"�,O5uB�����t�V�g�xL��ԓ�>72�����dL��֥���n+�s�?�'�ܼc�����Y��`8+>��*�d��LrJ.��_�fG�x�ЩT�q����ڽ��89%��g�B^ )�^S-HC��B>�7_�$�G>�ɶX'ҕ�>�QI |3�z4�޻N���d�!�����A%����,H�Q�
��̌ ���X�P�K $I��M�E�J��ŉ�J!�b����$mk��)�jʥBT���亐�W��Tlq+���@�$�*�xV@M��]�@%:=��H���)�f/щ�����=�Vx�+�q��!�XH/C¬�϶�YjzN�V@��6�ո��*��n��=4�E��W	.�|�2�X��p�m(���W��/��t��Kg�ڥ����^���;��.���r\=�?�C���/d+�8Mܾw܏V��؊�����ℹH|ee).�;_�ܧ���k�Pl���7��v�Q�M���eJ�^���6r����Z��O�h\��B���8�=�7��vl��vQ�(��wa�:�k8#��+���_�O~�U���)��^?�}��;�G��h�b���5�[M�ucc#^�eʽ�N����l��{�G�qA���N�9{:^��g�9�rF���d������ƣ[�`�F�\;�Ȥ��Ht	���K/ǵ�7��Kq�̙x�����O'm/���1=�Ŏ�[6.����V�r<��O�6��b<,(g��[qq���|+�#�� ��������a#��ބi|d>�Xk����8�i�u��:�Wfu�'X�˜��Ù�t��/����٩�C��8��$�s�	�8puV9�q�(q�Hώ4>�(e��3�ס�m[��"s�yy_=C��s:�/�,��6�M�#���(�s.>�6����ö�G�]S��p����w*YX��u��M[�[ӹF6_��͋sT#�{�F�Y6�Ҷ��+!gKu��Gk�Q&��} �ũ����N�?4i�Ի�����c��7�μ���~�y�#�_1�?mGt9��n��q�~��|���viY�#͡���)��M~!�6w�N;Vϣ7�]�� �T/|ϮL⳧��7���gO/��܇�?Kf}�~���%�$aB�'I�6��K2*��� v�	�#��+sf�u2h�R���df��!2?�`���#k�����p�o91�2�\D�(M���wr��d�Ӄ��� ʌ���e��"pc���M�^��g���"��|�O�U�lU���uF�*��u�}�O1����-�8�^ 
GҎv/��z��uzl�3������޻���.�s�;�OPkT�t�6P+yʨ�xa�3}���������g	��f,;IӒO�S�Y 1�[�d^�,��/�ܼd�d��|�7�hw*�����A��rq�
5m{Vo}�_���!G������_�:��Iҁo*Sq���Gi.���y]�u:�8�։��oǩ�g��Wnī7���>����^fqp|v�~�H���΍�Sg����ĕ�7���_�Ͼ���\[�	���il��W�3�y�1�![]ߌ�?���|�Ÿ|�����H�=�p���[�c`�/���A�������7���W��W����J��Cp���.����BuǙ�����ԥ+q���x�����ׯ��Gj������>��*t����N�&�x��������'?��_�7_�KW�G�����ѥ��3����$=z�[�&��'������'pB_�W^~%�_=��w�v4��ڵ�Z��Z���nl�;1�-D����|��gI���@9�BN��X�cӭ�,���b��wc��)�avV�ؠO]w� l�ά���o��9��Y�*�|'+��ɛ�F�	t��7[BI9H���ٯ,��,��dN.�S��k���T�C�&ҶC��a�ɝ|3�\���Rp�`Ud� ��Bl��q�'q.�X���ət
�C@|�u�L��Z�,�[��d �4���|��2��VI/���$zܫ+u� �阊΢ߤi4E�G����9�9���w���lx�Ƕ����X��v#�����F=���c>�a�b�kz�=Y�`�5q��T�-˿dIi��$M R�x�,��G���v�������3;��Vb�#�%$�'}���G�{��\(�yQ�f�݊�(��S?}�c�#3)i��!�e|;�b��HR����.��yӸe��X�p��g<���J�#ɐ�#�0\"+`�'�?����d�+C�E~�zVM��`��:C�@����Rǂ2m�Z���̑���%j�	8:uY�KGO�ý�H���~�({�(�'P��*$J2��,���|��F�c��()2y�Ѥ�.�I�ӻ(S���O@dI`C��6���+��2����ǦZ���d���ms� �xvK�[5 ��(�;I���h��!��%B�\�GE��^D*%���b�O%F��Q����
���0�%�f����8r���|�n>���%�gxx��8K�ц/��|!��~)�7�����ǒ����|oq{{w�=����8�ii�V�,N���/\�Sg/R�Z��g1��0Q��A#��q�΃x���s
��O>N]��k��/��֗��Z��0�����(>��$?ًѴ���ǫ��T\}��X߼�.^��6���鰟ߴ{��Q|��Vl�.�X������_z��\���Z�+g֣>��{s�Z|��a<>G�Z�\���z�
e��F�7�j���k�˱�b��^�O����a|��۱�ήݸv1n�|3VN��=t��n�;�W�.���iF�x�����Z�=�o{g
�ط�NL4�87��2Ay�u1�ɫ򲏠L��A�O?�� Y^�tF���@囹>ڊ�(�2�7�~^�g'���V1%�|>��yO)$s:��<���{�g���0����)��aU{��!'-g.��Gm����y۞�|�̩�c�,��6Z��
��,��t��n��5�m�e��\'�rC�8;�b)�K�	��	�<Łr�F'T���'�V�&�B�qk������7����!�,���9{(q�����"��� ��)���������
i���N˒&���7g��RqZκ�c+ˍEO1�<凣����-qɃ{�e���2;8�t��c�86��Z�V��3�Z/~�b/.-��V���~:mk+���$�?I�?��
 {��o<:����w㗷������3�b�rS \W�	
0�d4G1\�Y;Y��a�l�\a�i��K�.�5����i�+f�{�皂�~�#�[I
IqN���\�Bl���Y��*���_�M�IYH���̝%o�J��-��ϺP�cG!��u#�D!�I�;F[���484@a�c�ĉ28Qn	�k���0����U���?�X�J��i��9�ApVT�z�K!L��V%����І�^ɮ��lK(!�Ƹ�㥁��S9w�7������q� �'a��|�H�Q-?)8�OT**�t�+�PAe��b&����Iĥ������y�}�@�:�C8�VҒR4�~�^�W�rMNnV�H����(���8�����������ɽx�}��̧����1�z?Z�%�A������O�N���o\�O��bܼq1F�9+����T<�:���V����~���{���x��{����Ԍ�_{%~�?��A���_�����/��.�hԎ�����w��W���p�(�V}�37�/������R<��7�^�Ͻ�\��vۓV����?�O���=��q������|�~�Zt�{��Qz����ڥ�hNb{8���?;����Ń���Z݈�7/ǧ_��];8}�e��3yq�7^x.�^\��}�[�֝A��_�f|�G��|�k�/���Π�ߟ�S�Z߀���S����x��a���}���š>{y�ߧ��S��F�3��d���ȿ��>�W����d��Vx+��<ʁ��
<䬴1힯�cT0��/{�=F*��MVy�{`����c��7I>#Q�G����oqIv�G��5��i&�C�T{��!�\sF/Z]V̅�2��҆6+��(Z>�B������=To�3Xi�p�#K7��R�#�z�����g����'��ǸE�|�R}����y����GF�Y u A���(uC�)t���&���ns��V��v�>e 1�#�з��=m�NpMR��r�it�1�c�)O�2��%_`�>#�fE���Jq�v��
ڭ�A?�R��p3aŋ8�S?��"�C�i���[2���vX�	���m��uQ�O��~�h�E�9�`���^4��,��_����jG�����l��������?��OՉJ��GOPx#ek/~��N�����#�����b��]C��׬�h�E��q�g�lsvFO$eWƳ����6�b�4l2��JO��yR�g���3�R2��SP��1�N��μ2��!�}�GA�)d�&:ϘUea�oIye��?a&�Ʉ��[nF%��P��~�:2�Q���El[�Ѻ~H�(����(���J���F���`��|<e܈��Ld:|u��=�fg)�LQ���锺~F���Y����c��������o���S�
��;6ԷZr]y\�Q<hGv��2ǘ!�nK��[��_#W�V���R��y�<�#G��'y|d�<Q����ee�D9��X�@E��6��.?�����k��8�U1���\��&�o���回�����d��������)Jp��N���^���3?m�m����3���ί���O�����߉������Ώ����'_�Ͼr5j�C��z�v�\��vbx�������a�W����p�#Ԝ�k/=?�������V��g�̹F��,�?������W�W��.lٍe������g_�s+��~?.n���˛ѝ���A�1^������Ocw�sx�♕���d|��˱<ڏe��s�6Q��t�������;����$��C��˱�m��������b�2���n-V�8uj#�[���׾o?�?�7w��/ׯ���ſ��q}s-�8^����ȝ�b�1�;�}5n����[�/�}#t{m��� ��`v�w
arH�Ӏj�'8:���.�~J53:�Q䠇��S�*G��kahw�݌��N&�\�5<t��2"�a�:�<`ٜ���%�ҧ@�6f5�&�8u�^�>�p���;k5�9�!��8�9��o�«�����:��<�	v@�,�z@ݓ��l
�XP>0������V���:Ψ:�݃�����m�m-t�B�6{8���� X��㗏� ��Yη�	�с�:���\BB{?�4��C�ѿ�^Z��J���x������1<���Nqp���/��@���x�������7P}t���RZ��N�y�#������rw�k�X�c�>��6���;Oq�ԯ~�>H�Z8�Ȼz'?[� ���X�����kG�% u����ԋ,��8��S����F1���t���W�%�j�8ҭy�7�=�6,�fL�bm�E⮗�*r����`��=��V<�ҍ��gD^�s�1��%�.���g����>�N�i�@8��Qރ�ғ���Q�!7^���0�c�1�d��7������)B�ϫa?ꔪ
ŷ���M�:M����i\�!�3�u1�NG8d&G�GR	L�&.�R��(����P�B�1�Ys6�9�C	�����������۫F@����-�o/%���D���Ƒg��D�<��<���O#�C*ޥ�%���NG������]����M�j�=S)^�J�[�n�P9��>u$['�o�CI]���#�r=��D�prFcn�K������]��Ƈ*�	F	�Gz���o��낚�����W:��#y�'F'M@� ��M>逓|G^ʹxW��dtg����@r���_��E�a��z	���^*vbM��K�TL���Ȯ�U��^ $��ِW��G�sa'��R:U�9��(�1N��p7.4��k����s�Ў5�6�۱}�h� k��5�w��1@^�8!-�g7��+gb�v-��j'��Q�Ĥ�o!wߺ�4vj��.:3�z����2��3K��؇�Z|��V�֭����8��N�#�8���k/nƙ�g0½XCϭ�A���c������W?܎yw5庋!z��ٸtf#� �2�~f�lҏ�֓�Ӈo��>|{�%��B7,c_{ṸF����@5fc�Nt;��W�y�E;�6��N�\F�}�y�z\>�[��2N�����I������(4����!G��:�ש�a���ɨ���b|�}0�.�k�yYCo`�f��->�]�(������D��eҜB�]'q�����A-z�^ʃ�z�#/Q�}�&�)�4TTh�r(O�"S�qm}�A�&���GC� �/�}�\�p��1N�;�'��=�܇.u-�sk��٧�gRd�8�(M6��s�:��������x<&�t�uB�;w�S��������8���s�4u҉bp�oib���2'�q����~���m�.�j�>�dp������i�G�H�\ʡ��+ 3�=�q/5���hs��%/���o�Bwp;��d������1<:�Qk%vƭ������m��ǚ��F�zV'J}@�� (�/��� yډ��y�����u洣	/���K9�:©�5��2�F����6mR�U:�8�8�M`*z��3��vmK���� �ᤝ��Ϯ��o o��.xB�t��];�k�<�\.��	١0��9��;�V��q�j���)+�߁�=�3�Ng)�+�ZP&��Q�L�oe�|\ƽMM!˾+�ꍷ�1�sv"r�*� 垻俤�L�����i�T"�Ӆ��R�9Ňa޼�!0k��RA*!�r�ǿ�H%�}7�7$�V�7�#2�����L�ެ:~o*33:7�6\h�Q��x�8���Q�&��m-y�і�s�U��+m*:O��>�����yQ��I�e)`K�B?�+�6qhstSUX>kb~�X�l�Vn�Q���!mL/�^��m��2{���!GQ�{��>1�\g>R���,�F��d��(UKS��}o;АdJ3D��t��2���G����1G��U��8�A��y|�}de�|&:�gs������?��h}K8I�zM�̣�?��i-Ek�"�m�i<����p�I��I[.n�R���nnA0 �#��ً��2
�9�WLuPS���W���{��`?�Kk1i�g��Z���܆`0f{W1D�(���V�=�m��SWc�[}ײ���h��^�PJ��v�1|z+�������q����������A�o,� ��8f:���;��7��|��+?k_g��d�g�)gy���}�.���(�T����R�f��lq����kp��W�}�F�8�.|����,�3��+�ElQ�q]p�Tj+�k�r ��ʓWx>�
�@HY��d�|l�]�'��l���!L�k9g�z>n�e��������$�$��t�r ��G=�o��/,]*���� ���>x?��4%^��<��t�t}j�k\���_'�/Y��T���FܗR�c��C�Q��@_Bp߱\?ˡ�:�s����'�4J�=�\����-�3��P��3���q�b���j����֓���E�§�[�[>+6I��,� �A�_+�OhU�~�)�!y%�}�?U'�NX��u-�v��Tz-�BM�UsA"�S�2�#u��^����d�����q2,�$˳r�-w��D9<A敇�����2�n��l���Æg�}��V��a)�-�� {"3*x����P֞U�S@��B����d�^��M}o)�e��-��s�N{`Ϊ�t��ў��
�e$�m!��qa�;���]4+��R'(d�RQ4�`��+�wN��93&<�I�UJm+�i)��d>ϔ�p�/٘��*��H��3T#{��E  '�IDAT��{2�8ƙqq�j}y)g����Tf�k��t6���6��]>~QA���r]<���[�����z,���d�Mp4t��YW��r?��V�����nJW,o`��9�>����)��S�cm����ۏ?��׊^�l��ض��;�;z�N�GF�O����[��3ע�;-1z1J��c0�%~��>Y�^�zr�����~;��/�s�&6N��=�u�D%Ջ1u���ϣ��_�U�s/���q����Ё����B��ix�_��Hw�t���`{O�x���'�ja[>�a��I�m��gp�T�ZHY�X���:�aq6s�T�㟷N(�`>N擯�̏J��&kʯ�������ė�Y�1孧�.� Y�9��K�')��A�'۞Y3�nȈ�:��~�5d�EE��j��uYm:�Y$Na�f>˕ȏ�El���*�=(��7�:�<Id�~�X�aj��C�a5�+�I*N^�I��u�A���*#��U�T�"����,_��Qy����H{���`�𑤊,)�y.?�<�Q��b��`zQ^�\lY1<���(� Z�J�"mq�d/uG��m��z2�8*iU:
H$��̥�a�ė;��+�Siz���K�B����*�^TZ�׉��5˛P����UQ&��c|	\����B���+�b��;�'�"UE.���6�n���SG�*��Ƙѿ��c�O#�`�D�&*Wۣ;V3eI�m4�Dh�͕ʛ��3i����\#������i�qDqJt����ߵg�V'?dNgrN��D}z���Z�S1��W��X�Cj	K�\��m��h�v�<�no3:k�(�.#\/q*�~��.�⩥h�L��§���j�i���-]O~��]g��ҍ>�Γ��`;�˛1o���i�.�I9����:oK�F�����˖O]�y�44p� t�r0�sF���~K�V��ء�7~���^9���Fy�7�i�B�<��ߩ�J;$�v��[��g��ōW~0N��I��)y����"�aюҷ'�,��c
�y�q�]1�8�q��FP���?"Y��L�$��p�[G$JkJ�yUxO9""�̦�����ɴ�"��*�.d�4�	�����ŚOc|�e�|l]�Q�O>�-��A����:A����S��*��p���Э�8�=�-�m��ǂY��ԯ�y�H�2�{[�,,�Z�;�w�-�-"�ܿ_H'��B���	ԟ�2��3�Z~�������uH��/������?��p����)"��Q�)o}y�q���c�P��DO2�rm�b�Mg��<y�
'�?uY��-�'�rT`�u�'���Z)Ǭ�;�ˌ�wJ_ �hZbs��,�N�[�[~�m^���%�$�q5��?��Uҽ�W�O7��d�v",���i��1�c�B�p<�EЉZ��g��4�#E:����Lw:��׸�g�xe�q����E1��_.���=e͙#E�b<R�g}'����}�iS��d���4r���?�� �Ҹ׺�\_8���3����іfL�+џ���������h{'ec����8�ߊ:ej�31�4�0k@C��ڏ�^:���8��1�ac9���6`��CGgs�˝����q��-�A�O���|��/��U1x��u��D=��G��_:}%f-�(���)k�'}�,_�^�K�v�|���oEg�T\z��hm\�~/vqXur1�ɋ�&���;o�f�H���gc���j��4�����������3n�F��r��%
z��D����P�+ ���[ #�3�^�L�Oΐm�Y薹�2%�A�s��<\p���疓G�&3hd����aY�����$�g�[U�2Y���� �6Ӷf�L+(U<V�)��<�tX�e��g ��"+̒�2,JB�e5�Q^�Q:�J<��q����G9��x��u�Ծ���Cҹ4�`���]^J�Q�~<��U��8{_�&}���;'���t��'m�N� ŕ�4g>P�x�Zհy��^�H1��5 TI�)��+X��)�g�>ĉ�|��嵇�V�	��о#��N��.$=�K%H�R)-�h	o�E����ch�v�n?������k�oa�g�iȊ3s%�2���ۼ���2��yI0=g����RВ�5�-e͓ƌ����J�0�3�,�7,�R�\<���0���#�YI�d:�)'�N��8wj9��x|�]�W3����Z�q��ĳp��.�ԉZ��bz���$j�^4�v�7���Z�-�j+���Vj�V����H[���bV)�Y+F��[QB�Ub��1*!FDDDn����W������<�9�{���(Ne�۬��E?T�M=v(���T�k����)&�0�,b�f0Ʊ�W�w�!_�͖J{<��vW�Hn�h��7-ZR��x�����OJ1E���j��4&�_�<�k]��E�a+J�{�+M	�r�-�u��N<F�݂@Z�$�F0.~L˓�zt��d����}�,B��%��܆=J�2ۛL4ۀr��e���%ڿ�X��(���̓�'�R!7^M�V�??���,��ʌo6�<2&�P�_U����7��jIO�|�oUW�ߍ{B6����*2��37d�)��I��	����Xɶ������˫��Nak9R��M���}޸�ΏC�t�RM>���o���gќ[v���D��ʯ�<������a<U��T��	ZC����g/�=+j�SM�h�ƞ���t��5ܛ/��3Vߝ}�E
��--�u/�/�aKg�lM��w���B<�wJ;v0=.^F��Դ#zc�+5� (|bB�}sG����.�7�:JA�����(3���j�ݱ�'?�_�<z�o�B��ͨ��=Qw��乓�wF?X���18i��#4z:PSa��T��$%q���+���H0����'� ��/`�k�/�U�	.��Z
y�2��^�#�)�S?�Nt��q/T��OP��H�5�Qד����E��.�[��Ǉz�'V�	���I���aI���n��'�Mj���!ם=�h�`���k���Z�`��霙1M���7+�L�$!U+����	li!;}�,;�@/H7w�Z�&���Q˰�c�곑A% ��J�O��[�pm��r����CԴ��-�yR���a��I��i���ͷ}3&��u���2�~w�]�0\J�"�#�Ⱦ�M����u��tw��^5u����� K:6�ld2�����k D�����\vYNh�^����g!�޼U���ӟ2؟��Nſ�k'����P���E���0�������v]����
����\�L��=�C�&���lt�(,a�!��F�DF(\��WaCPu,��]��~s���Q<E�Fnj>����`��=Ѿ?��-�~�֮?a�e��t���	�ڝ:bB�m-̃�ڕ�{�g�ǚ�\��Y�Q1��˸��U'�#.�g��X�-ϩ2Jil������B�.�r�I�����]/�3$�P�K��Y�b7�c�-�Ȭ�̆N����85��%gP�H���ZwDô����q-��N��i��5u�{�)��>�������%J�6��-��\�`T�5ҥ�pJdu����]��P��W�D#�Xi�4�ϥ0���F���u�����1�z�X �7u��6NWpq4h��j��jC��mPݫ9�ѳ(�K�v�Wy)�~P�P�زp}����K4�PIqD�D&M�^HH9T��K��͖�@램�
W��C��}�4k7�'�禂�^�b�d�>�\�9F�k�C�ZE���O�8��r_��hR��F2p��={O�x�5Dȳlxe�y�D��:^2�L\�'���<��
� Q��M��@N�e�(	���7N��+��5�_g��-�T%cTa�k�v#�Z��ر�H�$�9ǉH�7��� ������e�(�s�n��N�e垡ٟ�P��u��n��E�m��{k�|'��
�ڙx��v����>Q��~�ߨ��ʧ��mq�Q�_��Jpyĭ
1W�>йd@cY��5��O�K,��n'O��p���4���~E�8��of��:@F�(�\S=�Wل��/i��jh��:]a�������ׇOD��[�=@9�K�a���-�\K��X��~�p�/}�qF��?+��#s�D.r�c>�{�G��G�M���Vi�܋��Ւx�d�=��]�[�I�+�~M�'1�W,�y�d�e�0	a�����.�U��߾k\ݞ�z�q�&I�=��k8���$���붮_���C���b�C�U��������(��h��mЎ���:����DQ-���RQ��K�oq�n�H�=Cs�+	Fb�b�7΄����v���s��:>
&_����|L��Q87��{I�4��*����a�s5��B��z��(C�5)_] �ߺ��v�
��<�(Z���]�G��L赨�&���'��:����=��cu������_Q��7�f���p�FX�j�g
nK�`�W8�_;"'�I뙁c�(F�O�᷷Z��!��ߝ��y�Q �����7�Rq�k?��̌��^��J�<�ۡ�x��J4�d>��Yv�n�~\ϵ:����tr<\�2F���O���B����1�3Ȅ"46s��`Q<4Mi��e<nB�P:>>$E�G���Ib� ա��>�|Zם��cIl��[O�l0h�O�4ݟy�̑�P�6��p@E�&8��I�@w�-�˷FZG$\3j�:@:�x?�ZNOR_�� !<�h[�b�H0J�]�)z�[��i+�x\�Gw�#<��Z�G���]��l�聎�R��d(�}��n���O���Lm���M����W�	��[�R�Z���ue#�F�y��7tn5��a�j�����c��,��M��y���%`�f�GG�P�m[���2mޜG�d��<��v�Ö�*��̕��JQH9!��������<Trh�/.5KM���(R�<�������ݮ�N�UCj��������<'˟�w���������O<������7���xmc���s���ܤ۲~��~��*V1cE��O�$�f��o�+=7��!�=��>�_��B�ۍ������3r�Y�g���H�I���o2@�6)���P�z��*���)ڃ;ϳ۴0d�liNq9�`�xdk����8ShъZ��Ք��eX����w|�Bxf�����Ƀ�d�\~�E�,��5��n��'��#�{��Ol���ڊ�srɧ�\H��c|�fb!i�V�O.:�-*y���y�&���@%��K�д���Dr�]t������E���[�>���7��*�?V�EWXS]'��Z�mٷ��Gܡ�d��6P�eV*O]<xk�)�Dՙ����	���Z���2�FuÐ������[��W����0���ddA�
�(�4g���#��b����.�L���zݪ��y�Y<�}�A�"�bc�(�AZ`}�a��4�U�b9���7.��|��J�lW��wn*ʪf�kj�PԂ��1����<2+s���[RT�xᡍ-?���7�f� �2���՘�01���SJsn�-ާ�D�+�+��^Rc1:3��!�' k�*Ǣ�����!�h�ԃ�6��F��+ՌO"�e�1��ۈI��o�����h��i0���dS��5�<j�2�6;�/���]�U�� d��]CE:�(�����C��H<�D���>.�,����q�t7.e�����(�a:tc)�6�����ZI��!���m�Q�NB���5_����W���I9��ǋ��Mx-���E7��?��L��U�"���*X���3J�X���թ�iFk�3Ճ��S�w,W�}��u��Y��u=̉�h%�("��00��E��5_J�)}��È+�-C��`��#�D���q\wu����qI��I�����3��X!&���]1R�mg���c�V�,v=����:j�T�"4��������}�Ө��x�Mv�(���62v��U��?=����ۈڢ�;�rGv�7�5]�;H��d�͌.W0u몫�!����.ô-������E]4��z
�d����S6�r$���k�=�4U�7�N��n���+��Ϳ�/-�̡�4��^]�"�sAH��Y!N;r"jJ�g��qYa�^Y�ށ� ���]����Dh&�MҲXQ���o8|.T��[��;=�R��9%���j���Fk�F�5�R��wV#��ط�G?�[ۨ�󭴻׋��6)I�^ċ��`��#!A#�~�=0��?l91
c�S�:+!�J'�j߇�C��Z3�G����f�dOI�T�[`S�ze�ւ ��(��p輻ꡚ�jXp�{Ża�?G)���)+��-�����O�y��/����'b�\�U�r�+�~�D柋��"�=����am��v_�9W�M)k�E{5�S��T��z�'���O���|k}�
M@����r=����1G�å��� egޚ)��ˌ}��;��U��a��m��T0�	���|�s��H���K+vkֻ���S�fY�"��ʣ�I��1��?^+�eg6��9�9�h�Վ`+�@�*����<���l�5�י��e�]%��N�����p2��Z:L:
����.{�b�C���=`v��dcg��$���ը#<l�ҡ��ܨs�����5����d2����#����ډ[��A�[�[����w����y;�����3Q6E��Y�ya�v*�U���ϟL
Uy�v�����QDV��9��~�{OÚ?�x��1�D����uqKG��OIҋJlՀ�z�ܹ�5t��s�,uīR�RmX*N��}F*g�q��m��3�D��I3P������[b�;�҄|��Ἆ��z/�#�`�mĔ�F���C�BH଼��+}^�s�֢�����7���օ_\Z�M�&X���U2�ѣ�m��C���V�6]q�������b���[,\���g��?��P+@F{��8}�<�MF5k�y^��nᕄ|f׸�z�7Ov�yItEO����Y;%�m-j8H?���.�S 10�6<�)l~n�W��%Y�zX�'�ƒnz� Ǔ�Я5��2��~O��H�3���k�Ӡ6� ���c���y'�#���?�q'+���Y?kM/5�h�ڝ���%ئ�}�`����縜��Աa[�^
Px���xh�C�O��~q�G��
,K��Z�~�UA�|9��E��;D�p.V7�h&u�Z��iݧt�]Lp�ž�v�Z�s	_iwcʭ���,�[�EB�z��5�4m۔����>�p��۲]���d�Mّ�[����AF�<�J��9�!��J�k�MڛI�����[+ŖJѩ��jc��]�9&�i�JGXV�6/:ȝ>X�[J h)�џ���5���IL?�nB=[��˂#��U�+��m��l��-�.? ���> �񤾭��!��Kd�a�x�콕e��m���w;��Dsĳ g�����JN�#����P�.Hq��c��,��9R����_/]jP�=#h��+lw-K�x��_E{��OYW�<P�m�"{P&��<T�V|�����A��u�����{3fH�D%��m~��%��X��s�n!Y�@���[i�/6�2-�=�|�Ilj��6q�^K��M�%�՛�S�b8\�E­���f.��.|�&��wT�җ����`��4u��3�n��rʞ݅��9K?�`w��{��	7 %�Y���5���
chOBaw�b��4�wr�1��e#�#����%̗�
~�u#�*Zlj��Ųd�Q���qLQ��K� �i�y���L�j�S���>��K̓33�����)-:D��dr�f߱�����|`�,����8�O��S�̟}yA��l��R�R�����6�D��۰�E��s-�1ì5V��ѓީ�ǓW�l8������I��A��F1�v��t���M�WV`s"��2ث؝�q�����,�'iA�t9�����9������J�|3`���^,��U�#.�?��.!Փ>�Z�9�K����
nA�]M(��I�uY�Z����_i{kC����$v9���A����fJ��e󬆟w�K�"f�"�l�r�*R��*uÌ-#=f��b��uĬj��O���)����G�֍��0�W�����}�X�T�ӳ����B�<Xļ�����|<��"a��;��o����rX9�9%�1Zi8���Ƨ�4�"TDU�B���Dw��{M)�F�ɓ�XMp=7h�3D@\[�\�F6�[���C�-�~2��Z.=;N܂��h�}��X�D=p���6�9����.�5��ns�E��蟟���8hca��T�=&0$�=�x+lǉR��芨���+5�3A?F��W�t6�}��[�iեk�Z�h�8*NF]`w�O���=���i{K�����ۋ2g�����<���L}p��n8PnLA�/"���;��w�`@�yD-�r��5�����20������5��Ѐ{��3��S��6��V;�U�D�kӑ��]���d(�
�3���wp�d����(�Y茘�edjX� @��8jɪ�����$��F�ρ�C3�/࣌�0������ʋ$D/c�܋����0Rk}��m��%���/��� S6@큸��n0)�"����)��s@�o�L���9�ÿ�>�9�ZQT��m��ر����,�|��j����n�]~���Y�Ҭ����S2�LF�/�̵����X�'��a��Bxo������D���9O,��+sn�?��䴝k&vZV�V�:S#L ��;�R�5�A9��dy���(+?�r��.�h�ps&��ő�
��|6�Dyt2gI�8S��O[V���`�ϛ�F��+A����D�'�Npm��Q #���)Z��0Od�hF��8
b�ʸ�PѳpF@@�M��Z,�Q���c��N��9?��L\U(���o���
<�h�97J�^����,-�j��8�RmX�؅����zDPoj���?�cv���|�B;fS\!ם��߬��+����:��	��,�:o��}�-.�1��t(9�	�)&���ں鸆��G�
A����.�߄�3�/$\�ZY�.jSr`���OFƉ�����g�r]d��Eڡ�o]�a(&�Tzdj�7�^U�:-�Akk9�b;*#*��iL��/>��yۧ������o.I��(�Y�7����$�vd�#��v+H���+1,cy�K��� ��X����j�d��Zљ���~���#L�����s����Z�D%{A��Y��s�7�����da���y�I�j	�E&�Kq�L1��7+�������LO������?'��j�EϮh��x�2�O�hj�i���_PK   m��V��'�W  >     jsons/user_defined.json���n�0�_%����lU�dhU��TE?&�DljC�(��{��ȐV��{Χc�sBͱ�(A������Ҳ@���)�aA0�&��z�C������{�r��,���X�i#w�A�^��X�P�R�y�BF��܏"�����OEGy,�\�����Ic[��a%]nU݌/ٞT~#�z�Z�.JNH���ru��M�D!ǜDa ��nc�.Ą1㕴Z}�A����*�'h�����'���<JY�y@9�rw:�0���Vi&{��t>���eZ�[��ψS��OɄ�9�ӷ��`z?K��v�G_Ɩ��6u0����QC��b�F��>ݶ�PK
   m��V!je�  #�                   cirkitFile.jsonPK
   V��V�O.2 �' /             '  images/7863607e-9197-4466-b19d-a9b84c893c9f.pngPK
   m��V��'�W  >               �. jsons/user_defined.jsonPK      �   20   